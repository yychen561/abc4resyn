// Benchmark "i10" written by ABC on Sun Jan 19 15:24:39 2025

module i10 ( 
    \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) , \V10(0) ,
    \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) , \V248(0) ,
    \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) , \V66(0) ,
    \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) , \V45(0) ,
    \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) , \V34(0) ,
    \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) , \V293(0) ,
    \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) , \V275(0) ,
    \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) , \V257(4) ,
    \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) , \V149(3) ,
    \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) , \V165(6) ,
    \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) , \V169(0) ,
    \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) , \V165(3) ,
    \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) , \V288(4) ,
    \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) , \V229(3) ,
    \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) , \V223(3) ,
    \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) , \V189(3) ,
    \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) , \V183(3) ,
    \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) , \V239(2) ,
    \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) , \V234(1) ,
    \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) , \V199(0) ,
    \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) , \V257(0) ,
    \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) , \V32(10) ,
    \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) , \V84(2) ,
    \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) , \V14(0) ,
    \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) , \V213(1) ,
    \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) , \V8(0) ,
    \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) ,
    \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) ,
    \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) ,
    \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) ,
    \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) ,
    \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) ,
    \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) ,
    \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) ,
    \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) ,
    \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) ,
    \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) ,
    \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) ,
    \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) ,
    \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) ,
    \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) ,
    \V78(0) , \V94(0) , \V94(1) ,
    \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) ,
    \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) ,
    V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546,
    V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) ,
    \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587,
    \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630,
    \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781,
    V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) ,
    \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) ,
    \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) ,
    \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) ,
    \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) ,
    \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) ,
    \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378,
    V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) ,
    \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) ,
    \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539,
    \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) ,
    \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) ,
    \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) ,
    V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) ,
    \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) ,
    \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) ,
    \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832,
    \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) ,
    \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) ,
    \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) ,
    \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) ,
    \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653,
    V654, V655, V656, V1370, V1371, V1372, V1373, V1374  );
  input  \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) ,
    \V10(0) , \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) ,
    \V248(0) , \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) ,
    \V66(0) , \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) ,
    \V45(0) , \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) ,
    \V34(0) , \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) ,
    \V293(0) , \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) ,
    \V275(0) , \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) ,
    \V257(4) , \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) ,
    \V149(3) , \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) ,
    \V165(6) , \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) ,
    \V169(0) , \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) ,
    \V165(3) , \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) ,
    \V288(4) , \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) ,
    \V229(3) , \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) ,
    \V223(3) , \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) ,
    \V189(3) , \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) ,
    \V183(3) , \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) ,
    \V239(2) , \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) ,
    \V234(1) , \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) ,
    \V199(0) , \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) ,
    \V257(0) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) ,
    \V32(10) , \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) ,
    \V84(2) , \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) ,
    \V14(0) , \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) ,
    \V213(1) , \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) ,
    \V8(0) , \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) ,
    \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) ,
    \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) ,
    \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) ,
    \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) ,
    \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) ,
    \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) ,
    \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) ,
    \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) ,
    \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) ,
    \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) ,
    \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) ,
    \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) ,
    \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) ,
    \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) ,
    \V78(0) , \V94(0) , \V94(1) ;
  output \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) ,
    \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) ,
    V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546,
    V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) ,
    \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587,
    \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630,
    \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781,
    V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) ,
    \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) ,
    \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) ,
    \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) ,
    \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) ,
    \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) ,
    \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378,
    V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) ,
    \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) ,
    \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539,
    \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) ,
    \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) ,
    \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) ,
    V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) ,
    \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) ,
    \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) ,
    \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832,
    \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) ,
    \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) ,
    \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) ,
    \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) ,
    \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653,
    V654, V655, V656, V1370, V1371, V1372, V1373, V1374;
  wire new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1279,
    new_n1280, new_n1281, new_n1289, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1383, new_n1384,
    new_n1385, new_n1386, new_n1387, new_n1388, new_n1389, new_n1390,
    new_n1391, new_n1392, new_n1393, new_n1394, new_n1395, new_n1396,
    new_n1397, new_n1398, new_n1399, new_n1400, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1408, new_n1409,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1477, new_n1479, new_n1480,
    new_n1481, new_n1482, new_n1483, new_n1484, new_n1485, new_n1486,
    new_n1487, new_n1488, new_n1489, new_n1490, new_n1491, new_n1492,
    new_n1493, new_n1494, new_n1495, new_n1496, new_n1497, new_n1498,
    new_n1499, new_n1500, new_n1501, new_n1502, new_n1503, new_n1504,
    new_n1505, new_n1506, new_n1507, new_n1508, new_n1509, new_n1510,
    new_n1511, new_n1512, new_n1513, new_n1514, new_n1515, new_n1516,
    new_n1517, new_n1518, new_n1519, new_n1520, new_n1521, new_n1522,
    new_n1523, new_n1524, new_n1525, new_n1526, new_n1527, new_n1528,
    new_n1529, new_n1530, new_n1531, new_n1532, new_n1533, new_n1534,
    new_n1535, new_n1536, new_n1537, new_n1538, new_n1539, new_n1540,
    new_n1541, new_n1542, new_n1543, new_n1544, new_n1545, new_n1546,
    new_n1547, new_n1548, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1554, new_n1555, new_n1556, new_n1557, new_n1558,
    new_n1559, new_n1560, new_n1561, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1566, new_n1567, new_n1568, new_n1569, new_n1570,
    new_n1571, new_n1572, new_n1573, new_n1574, new_n1575, new_n1576,
    new_n1577, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1584, new_n1585, new_n1586, new_n1587, new_n1588,
    new_n1589, new_n1590, new_n1591, new_n1592, new_n1593, new_n1594,
    new_n1595, new_n1596, new_n1597, new_n1598, new_n1599, new_n1600,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613,
    new_n1614, new_n1615, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1633, new_n1635, new_n1636,
    new_n1637, new_n1638, new_n1639, new_n1640, new_n1642, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654, new_n1655,
    new_n1661, new_n1662, new_n1663, new_n1664, new_n1665, new_n1666,
    new_n1667, new_n1668, new_n1669, new_n1670, new_n1671, new_n1672,
    new_n1673, new_n1674, new_n1675, new_n1676, new_n1677, new_n1678,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1727, new_n1728, new_n1729, new_n1730, new_n1731, new_n1732,
    new_n1733, new_n1734, new_n1735, new_n1736, new_n1737, new_n1738,
    new_n1739, new_n1740, new_n1741, new_n1742, new_n1743, new_n1744,
    new_n1745, new_n1746, new_n1747, new_n1748, new_n1749, new_n1750,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1805, new_n1806, new_n1807, new_n1808, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1816,
    new_n1817, new_n1818, new_n1819, new_n1820, new_n1821, new_n1822,
    new_n1823, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1829, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1887, new_n1888,
    new_n1889, new_n1890, new_n1891, new_n1892, new_n1893, new_n1894,
    new_n1895, new_n1896, new_n1897, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1955, new_n1956, new_n1957, new_n1958,
    new_n1959, new_n1960, new_n1961, new_n1962, new_n1963, new_n1964,
    new_n1965, new_n1966, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1990,
    new_n1991, new_n1992, new_n1993, new_n1994, new_n1995, new_n1996,
    new_n1997, new_n1998, new_n1999, new_n2000, new_n2001, new_n2003,
    new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015,
    new_n2016, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021,
    new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027,
    new_n2028, new_n2029, new_n2030, new_n2031, new_n2032, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039,
    new_n2040, new_n2041, new_n2042, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089,
    new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2139, new_n2140,
    new_n2141, new_n2142, new_n2143, new_n2145, new_n2146, new_n2147,
    new_n2148, new_n2149, new_n2150, new_n2151, new_n2152, new_n2153,
    new_n2154, new_n2155, new_n2156, new_n2157, new_n2158, new_n2159,
    new_n2161, new_n2163, new_n2164, new_n2165, new_n2166, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2178, new_n2179, new_n2180, new_n2181, new_n2183,
    new_n2184, new_n2185, new_n2186, new_n2187, new_n2188, new_n2189,
    new_n2190, new_n2191, new_n2192, new_n2193, new_n2195, new_n2196,
    new_n2197, new_n2199, new_n2200, new_n2202, new_n2203, new_n2204,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2259, new_n2261,
    new_n2262, new_n2263, new_n2264, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2329, new_n2330, new_n2331, new_n2332,
    new_n2333, new_n2334, new_n2335, new_n2336, new_n2337, new_n2338,
    new_n2339, new_n2342, new_n2343, new_n2344, new_n2346, new_n2347,
    new_n2348, new_n2349, new_n2350, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2375,
    new_n2376, new_n2377, new_n2378, new_n2379, new_n2380, new_n2381,
    new_n2382, new_n2383, new_n2384, new_n2385, new_n2386, new_n2387,
    new_n2388, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2449, new_n2450, new_n2451, new_n2452,
    new_n2453, new_n2455, new_n2456, new_n2457, new_n2458, new_n2459,
    new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2481,
    new_n2483, new_n2484, new_n2485, new_n2486, new_n2487, new_n2488,
    new_n2489, new_n2490, new_n2491, new_n2492, new_n2493, new_n2494,
    new_n2495, new_n2496, new_n2498, new_n2499, new_n2500, new_n2502,
    new_n2503, new_n2504, new_n2505, new_n2507, new_n2508, new_n2509,
    new_n2510, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2525, new_n2527,
    new_n2528, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2542,
    new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2548,
    new_n2550, new_n2551, new_n2552, new_n2553, new_n2554, new_n2555,
    new_n2556, new_n2558, new_n2559, new_n2561, new_n2562, new_n2563,
    new_n2564, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2592, new_n2593, new_n2594, new_n2595, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2602, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2614, new_n2615, new_n2616,
    new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2622,
    new_n2624, new_n2626, new_n2627, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2645,
    new_n2646, new_n2648, new_n2649, new_n2650, new_n2651, new_n2652,
    new_n2653, new_n2655, new_n2656, new_n2657, new_n2658, new_n2659,
    new_n2660, new_n2661, new_n2662, new_n2663, new_n2664, new_n2665,
    new_n2666, new_n2667, new_n2668, new_n2669, new_n2670, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703,
    new_n2704, new_n2705, new_n2706, new_n2707, new_n2708, new_n2709,
    new_n2710, new_n2711, new_n2712, new_n2713, new_n2714, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2757, new_n2758, new_n2759, new_n2760,
    new_n2761, new_n2762, new_n2763, new_n2764, new_n2765, new_n2766,
    new_n2767, new_n2768, new_n2769, new_n2770, new_n2771, new_n2772,
    new_n2773, new_n2774, new_n2776, new_n2777, new_n2778, new_n2779,
    new_n2780, new_n2781, new_n2782, new_n2783, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2812, new_n2813, new_n2814,
    new_n2815, new_n2816, new_n2817, new_n2818, new_n2819, new_n2820,
    new_n2821, new_n2822, new_n2823, new_n2825, new_n2826, new_n2827,
    new_n2828, new_n2829, new_n2830, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2842, new_n2843, new_n2844, new_n2845, new_n2846, new_n2847,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2858, new_n2859, new_n2860, new_n2861,
    new_n2862, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2872, new_n2873, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2880, new_n2881, new_n2882, new_n2883,
    new_n2884, new_n2885, new_n2886, new_n2887, new_n2888, new_n2889,
    new_n2890, new_n2891, new_n2892, new_n2893, new_n2894, new_n2895,
    new_n2896, new_n2897, new_n2898, new_n2899, new_n2900, new_n2901,
    new_n2902, new_n2903, new_n2904, new_n2905, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2930, new_n2931, new_n2932, new_n2933, new_n2934, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2942, new_n2943,
    new_n2944, new_n2945, new_n2946, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2968, new_n2969, new_n2971, new_n2972,
    new_n2974, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2983, new_n2984, new_n2985, new_n2986, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2993, new_n2994, new_n2995,
    new_n2996, new_n2998, new_n2999, new_n3000, new_n3001, new_n3003,
    new_n3004, new_n3005, new_n3006, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3013, new_n3014, new_n3015, new_n3016, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3023, new_n3024, new_n3025,
    new_n3026, new_n3028, new_n3029, new_n3030, new_n3031, new_n3033,
    new_n3034, new_n3035, new_n3036, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3043, new_n3044, new_n3045, new_n3046, new_n3048,
    new_n3049, new_n3051, new_n3052, new_n3053, new_n3054, new_n3056,
    new_n3057, new_n3058, new_n3060, new_n3061, new_n3063, new_n3064,
    new_n3066, new_n3067, new_n3069, new_n3071, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3083, new_n3084, new_n3085, new_n3086, new_n3087,
    new_n3088, new_n3089, new_n3090, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3102, new_n3103, new_n3104, new_n3105, new_n3106, new_n3107,
    new_n3108, new_n3109, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3117, new_n3118, new_n3119, new_n3120, new_n3122,
    new_n3123, new_n3124, new_n3125, new_n3127, new_n3128, new_n3129,
    new_n3131, new_n3132, new_n3133, new_n3135, new_n3136, new_n3138,
    new_n3139, new_n3141, new_n3142, new_n3143, new_n3144, new_n3146,
    new_n3147, new_n3148, new_n3150, new_n3151, new_n3152, new_n3154,
    new_n3155;
  assign new_n482 = \V149(4)  & ~\V149(0) ;
  assign new_n483 = \V149(1)  & new_n482;
  assign new_n484 = \V149(2)  & new_n483;
  assign new_n485 = ~\V149(3)  & new_n484;
  assign new_n486 = ~\V149(0)  & ~\V149(2) ;
  assign new_n487 = ~\V149(1)  & new_n486;
  assign new_n488 = \V149(1)  & ~\V149(2) ;
  assign new_n489 = ~\V149(0)  & new_n488;
  assign new_n490 = \V149(7)  & \V149(5) ;
  assign new_n491 = ~\V149(3)  & new_n490;
  assign new_n492 = new_n489 & new_n491;
  assign new_n493 = \V149(4)  & new_n492;
  assign new_n494 = \V149(6)  & new_n493;
  assign new_n495 = ~\V149(7)  & \V149(5) ;
  assign new_n496 = ~\V149(3)  & new_n495;
  assign new_n497 = new_n489 & new_n496;
  assign new_n498 = \V149(4)  & new_n497;
  assign new_n499 = \V149(6)  & new_n498;
  assign new_n500 = ~new_n494 & ~new_n499;
  assign \V802(0)  = \V52(0)  | \V51(0) ;
  assign new_n502 = ~\V55(0)  & ~new_n500;
  assign new_n503 = ~\V802(0)  & new_n502;
  assign new_n504 = ~new_n485 & ~new_n487;
  assign new_n505 = ~new_n503 & new_n504;
  assign new_n506 = \V70(0)  & ~\V165(5) ;
  assign new_n507 = \V165(3)  & new_n506;
  assign new_n508 = ~\V165(4)  & new_n507;
  assign new_n509 = ~\V165(6)  & new_n508;
  assign new_n510 = \V169(0)  & ~new_n505;
  assign new_n511 = ~\V291(0)  & new_n510;
  assign new_n512 = ~new_n509 & new_n511;
  assign V763 = ~\V292(0)  & new_n512;
  assign new_n514 = \V70(0)  & \V165(7) ;
  assign new_n515 = \V261(0)  & new_n514;
  assign new_n516 = \V165(5)  & new_n515;
  assign new_n517 = \V165(3)  & new_n516;
  assign new_n518 = \V165(4)  & new_n517;
  assign new_n519 = \V165(6)  & new_n518;
  assign new_n520 = \V165(0)  & new_n519;
  assign new_n521 = \V165(1)  & new_n520;
  assign new_n522 = \V165(2)  & new_n521;
  assign new_n523 = V763 & new_n522;
  assign new_n524 = \V165(6)  & \V165(7) ;
  assign new_n525 = \V165(5)  & new_n524;
  assign new_n526 = \V165(3)  & new_n525;
  assign new_n527 = \V165(4)  & new_n526;
  assign new_n528 = \V261(0)  & new_n527;
  assign new_n529 = ~\V204(0)  & new_n528;
  assign new_n530 = \V165(0)  & new_n529;
  assign new_n531 = \V165(1)  & new_n530;
  assign new_n532 = \V165(2)  & new_n531;
  assign new_n533 = ~new_n523 & ~new_n532;
  assign new_n534 = ~\V262(0)  & new_n533;
  assign new_n535 = \V149(2)  & \V149(3) ;
  assign new_n536 = \V149(1)  & new_n535;
  assign new_n537 = ~\V149(0)  & new_n536;
  assign new_n538 = ~\V174(0)  & new_n485;
  assign new_n539 = \V277(0)  & new_n538;
  assign new_n540 = \V278(0)  & ~new_n539;
  assign new_n541 = new_n537 & ~new_n540;
  assign new_n542 = ~\V59(0)  & new_n541;
  assign new_n543 = ~\V149(1)  & \V149(2) ;
  assign new_n544 = ~\V149(0)  & new_n543;
  assign new_n545 = ~new_n487 & ~new_n544;
  assign new_n546 = ~\V149(4)  & ~\V149(0) ;
  assign new_n547 = \V149(1)  & new_n546;
  assign new_n548 = \V149(2)  & new_n547;
  assign new_n549 = ~\V149(3)  & new_n548;
  assign new_n550 = ~new_n538 & new_n545;
  assign new_n551 = ~new_n549 & new_n550;
  assign new_n552 = ~\V174(0)  & ~new_n551;
  assign new_n553 = new_n537 & new_n540;
  assign new_n554 = ~\V59(0)  & ~\V60(0) ;
  assign new_n555 = new_n541 & ~new_n554;
  assign new_n556 = ~new_n552 & ~new_n553;
  assign new_n557 = ~new_n555 & new_n556;
  assign new_n558 = \V257(7)  & ~new_n534;
  assign new_n559 = ~new_n542 & new_n558;
  assign new_n560 = new_n557 & new_n559;
  assign new_n561 = ~\V59(0)  & \V149(4) ;
  assign new_n562 = ~new_n540 & new_n561;
  assign new_n563 = new_n537 & new_n562;
  assign new_n564 = new_n534 & new_n563;
  assign new_n565 = new_n557 & new_n564;
  assign new_n566 = ~new_n537 & ~new_n538;
  assign new_n567 = ~new_n549 & new_n566;
  assign new_n568 = \V234(0)  & ~new_n545;
  assign new_n569 = new_n567 & new_n568;
  assign new_n570 = \V194(0)  & new_n545;
  assign new_n571 = ~new_n567 & new_n570;
  assign new_n572 = ~new_n569 & ~new_n571;
  assign new_n573 = new_n534 & ~new_n572;
  assign new_n574 = ~new_n542 & new_n573;
  assign new_n575 = ~new_n557 & new_n574;
  assign new_n576 = ~new_n560 & ~new_n565;
  assign new_n577 = ~new_n575 & new_n576;
  assign new_n578 = V763 & new_n534;
  assign new_n579 = ~new_n577 & ~new_n578;
  assign new_n580 = ~new_n578 & new_n579;
  assign new_n581 = ~\V56(0)  & ~\V59(0) ;
  assign new_n582 = ~\V60(0)  & new_n581;
  assign new_n583 = V763 & ~new_n582;
  assign new_n584 = \V32(2)  & new_n583;
  assign new_n585 = \V32(5)  & ~new_n583;
  assign new_n586 = ~new_n583 & new_n585;
  assign new_n587 = ~new_n584 & ~new_n586;
  assign new_n588 = new_n578 & ~new_n587;
  assign new_n589 = new_n578 & new_n588;
  assign new_n590 = ~new_n580 & ~new_n589;
  assign new_n591 = \V149(3)  & new_n544;
  assign new_n592 = ~new_n538 & ~new_n591;
  assign new_n593 = \V60(0)  & ~new_n592;
  assign new_n594 = \V149(7)  & ~\V149(5) ;
  assign new_n595 = ~\V149(3)  & new_n594;
  assign new_n596 = new_n489 & new_n595;
  assign new_n597 = \V149(4)  & new_n596;
  assign new_n598 = \V149(6)  & new_n597;
  assign new_n599 = ~\V174(0)  & new_n487;
  assign new_n600 = ~\V149(4)  & ~\V149(3) ;
  assign new_n601 = new_n599 & new_n600;
  assign new_n602 = \V149(5)  & new_n601;
  assign new_n603 = \V88(2)  & new_n602;
  assign new_n604 = ~\V88(3)  & new_n603;
  assign new_n605 = ~\V88(2)  & new_n602;
  assign new_n606 = ~\V88(3)  & new_n605;
  assign V707 = ~\V149(3)  & new_n599;
  assign new_n608 = ~\V149(5)  & ~\V149(4) ;
  assign new_n609 = V707 & new_n608;
  assign new_n610 = \V88(2)  & new_n609;
  assign new_n611 = ~\V88(3)  & new_n610;
  assign new_n612 = \V149(5)  & V707;
  assign new_n613 = \V149(4)  & new_n612;
  assign new_n614 = ~\V149(5)  & V707;
  assign new_n615 = \V149(4)  & new_n614;
  assign new_n616 = ~\V88(2)  & new_n609;
  assign new_n617 = \V88(3)  & new_n616;
  assign new_n618 = \V88(3)  & new_n610;
  assign new_n619 = \V88(3)  & new_n605;
  assign new_n620 = ~new_n611 & ~new_n613;
  assign new_n621 = ~new_n604 & ~new_n606;
  assign new_n622 = new_n620 & new_n621;
  assign new_n623 = ~new_n618 & ~new_n619;
  assign new_n624 = ~new_n615 & ~new_n617;
  assign new_n625 = new_n623 & new_n624;
  assign new_n626 = new_n622 & new_n625;
  assign new_n627 = \V169(1)  & ~new_n545;
  assign new_n628 = ~new_n626 & new_n627;
  assign new_n629 = \V60(0)  & new_n628;
  assign new_n630 = \V149(3)  & new_n599;
  assign new_n631 = new_n627 & new_n630;
  assign new_n632 = \V60(0)  & new_n631;
  assign new_n633 = \V56(0)  & new_n631;
  assign new_n634 = \V56(0)  & new_n628;
  assign new_n635 = ~new_n633 & ~new_n634;
  assign new_n636 = ~new_n629 & ~new_n632;
  assign new_n637 = new_n635 & new_n636;
  assign new_n638 = new_n538 & ~new_n540;
  assign new_n639 = ~\V149(5)  & ~\V149(3) ;
  assign new_n640 = new_n544 & new_n639;
  assign new_n641 = \V149(4)  & new_n640;
  assign new_n642 = ~\V149(4)  & new_n640;
  assign new_n643 = \V149(5)  & ~\V149(3) ;
  assign new_n644 = new_n544 & new_n643;
  assign new_n645 = ~\V149(4)  & new_n644;
  assign new_n646 = ~new_n641 & ~new_n642;
  assign new_n647 = ~new_n645 & new_n646;
  assign new_n648 = ~new_n591 & new_n626;
  assign new_n649 = ~new_n638 & new_n647;
  assign new_n650 = ~new_n630 & new_n649;
  assign new_n651 = new_n648 & new_n650;
  assign new_n652 = ~\V56(0)  & ~\V53(0) ;
  assign new_n653 = ~\V57(0)  & new_n652;
  assign new_n654 = new_n637 & ~new_n651;
  assign new_n655 = ~new_n653 & new_n654;
  assign new_n656 = new_n534 & ~new_n549;
  assign new_n657 = ~new_n537 & new_n656;
  assign new_n658 = \V53(0)  & new_n657;
  assign new_n659 = ~\V56(0)  & new_n658;
  assign new_n660 = ~new_n598 & ~new_n655;
  assign new_n661 = ~new_n659 & new_n660;
  assign new_n662 = ~new_n593 & ~new_n661;
  assign new_n663 = ~new_n590 & ~new_n662;
  assign new_n664 = new_n661 & new_n663;
  assign new_n665 = \V78(4)  & new_n662;
  assign new_n666 = ~new_n661 & new_n665;
  assign \V321(2)  = ~new_n664 & ~new_n666;
  assign new_n668 = ~\V149(7)  & ~\V149(5) ;
  assign new_n669 = \V149(3)  & new_n668;
  assign new_n670 = new_n489 & new_n669;
  assign new_n671 = ~\V149(4)  & new_n670;
  assign new_n672 = ~\V149(6)  & new_n671;
  assign new_n673 = ~\V802(0)  & new_n672;
  assign new_n674 = new_n534 & ~new_n673;
  assign new_n675 = ~\V288(0)  & \V288(1) ;
  assign new_n676 = ~\V288(2)  & \V288(3) ;
  assign new_n677 = ~\V288(4)  & \V288(5) ;
  assign new_n678 = ~\V288(6)  & \V288(7) ;
  assign new_n679 = new_n677 & new_n678;
  assign new_n680 = ~new_n677 & ~new_n678;
  assign new_n681 = ~new_n679 & ~new_n680;
  assign new_n682 = new_n676 & new_n681;
  assign new_n683 = ~new_n676 & ~new_n681;
  assign new_n684 = ~new_n682 & ~new_n683;
  assign new_n685 = new_n675 & new_n684;
  assign new_n686 = ~new_n675 & ~new_n684;
  assign new_n687 = ~new_n685 & ~new_n686;
  assign new_n688 = new_n675 & ~new_n687;
  assign new_n689 = new_n675 & new_n688;
  assign new_n690 = \V288(0)  & ~\V288(1) ;
  assign new_n691 = ~new_n687 & new_n690;
  assign new_n692 = new_n690 & new_n691;
  assign new_n693 = ~new_n687 & ~new_n690;
  assign new_n694 = ~new_n690 & new_n693;
  assign new_n695 = ~new_n692 & ~new_n694;
  assign new_n696 = ~new_n675 & new_n695;
  assign new_n697 = ~new_n675 & new_n696;
  assign new_n698 = ~new_n689 & ~new_n697;
  assign new_n699 = \V223(3)  & ~new_n545;
  assign new_n700 = new_n567 & new_n699;
  assign new_n701 = \V183(3)  & new_n545;
  assign new_n702 = ~new_n567 & new_n701;
  assign new_n703 = ~new_n700 & ~new_n702;
  assign new_n704 = ~new_n557 & ~new_n578;
  assign new_n705 = ~new_n703 & new_n704;
  assign new_n706 = new_n534 & new_n705;
  assign new_n707 = ~new_n542 & new_n706;
  assign new_n708 = ~new_n578 & new_n707;
  assign new_n709 = ~new_n662 & new_n708;
  assign new_n710 = new_n661 & new_n709;
  assign new_n711 = \V32(3)  & new_n662;
  assign new_n712 = ~new_n661 & new_n711;
  assign \V1213(3)  = new_n710 | new_n712;
  assign new_n714 = ~new_n698 & ~\V1213(3) ;
  assign new_n715 = new_n698 & \V1213(3) ;
  assign new_n716 = ~new_n714 & ~new_n715;
  assign new_n717 = \V288(2)  & ~\V288(3) ;
  assign new_n718 = \V288(4)  & ~\V288(5) ;
  assign new_n719 = \V288(6)  & ~\V288(7) ;
  assign new_n720 = ~new_n678 & ~new_n719;
  assign new_n721 = new_n718 & ~new_n720;
  assign new_n722 = ~new_n718 & new_n720;
  assign new_n723 = ~new_n721 & ~new_n722;
  assign new_n724 = new_n677 & ~new_n678;
  assign new_n725 = ~new_n723 & ~new_n724;
  assign new_n726 = new_n723 & new_n724;
  assign new_n727 = ~new_n725 & ~new_n726;
  assign new_n728 = new_n717 & new_n727;
  assign new_n729 = ~new_n717 & ~new_n727;
  assign new_n730 = ~new_n728 & ~new_n729;
  assign new_n731 = new_n676 & ~new_n681;
  assign new_n732 = ~new_n730 & ~new_n731;
  assign new_n733 = new_n730 & new_n731;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign new_n735 = new_n690 & ~new_n734;
  assign new_n736 = new_n675 & ~new_n684;
  assign new_n737 = new_n690 & new_n736;
  assign new_n738 = ~new_n734 & new_n736;
  assign new_n739 = ~new_n735 & ~new_n737;
  assign new_n740 = ~new_n738 & new_n739;
  assign new_n741 = \V288(0)  & \V288(1) ;
  assign new_n742 = new_n717 & ~new_n727;
  assign new_n743 = new_n717 & new_n731;
  assign new_n744 = ~new_n727 & new_n731;
  assign new_n745 = ~new_n742 & ~new_n743;
  assign new_n746 = ~new_n744 & new_n745;
  assign new_n747 = \V288(2)  & \V288(3) ;
  assign new_n748 = new_n718 & new_n720;
  assign new_n749 = new_n718 & new_n724;
  assign new_n750 = new_n720 & new_n724;
  assign new_n751 = ~new_n748 & ~new_n749;
  assign new_n752 = ~new_n750 & new_n751;
  assign new_n753 = \V288(4)  & \V288(5) ;
  assign new_n754 = ~\V288(6)  & ~\V288(7) ;
  assign new_n755 = new_n753 & ~new_n754;
  assign new_n756 = ~new_n753 & new_n754;
  assign new_n757 = ~new_n755 & ~new_n756;
  assign new_n758 = ~new_n752 & new_n757;
  assign new_n759 = new_n752 & ~new_n757;
  assign new_n760 = ~new_n758 & ~new_n759;
  assign new_n761 = new_n747 & new_n760;
  assign new_n762 = ~new_n747 & ~new_n760;
  assign new_n763 = ~new_n761 & ~new_n762;
  assign new_n764 = ~new_n746 & new_n763;
  assign new_n765 = new_n746 & ~new_n763;
  assign new_n766 = ~new_n764 & ~new_n765;
  assign new_n767 = new_n741 & new_n766;
  assign new_n768 = ~new_n741 & ~new_n766;
  assign new_n769 = ~new_n767 & ~new_n768;
  assign new_n770 = ~new_n740 & new_n769;
  assign new_n771 = new_n740 & ~new_n769;
  assign new_n772 = ~new_n770 & ~new_n771;
  assign new_n773 = new_n675 & ~new_n772;
  assign new_n774 = new_n675 & new_n773;
  assign new_n775 = new_n690 & ~new_n772;
  assign new_n776 = new_n690 & new_n775;
  assign new_n777 = new_n690 & new_n734;
  assign new_n778 = ~new_n690 & ~new_n734;
  assign new_n779 = ~new_n777 & ~new_n778;
  assign new_n780 = ~new_n736 & ~new_n779;
  assign new_n781 = new_n736 & new_n779;
  assign new_n782 = ~new_n780 & ~new_n781;
  assign new_n783 = new_n687 & new_n782;
  assign new_n784 = ~new_n772 & ~new_n783;
  assign new_n785 = new_n772 & new_n783;
  assign new_n786 = ~new_n784 & ~new_n785;
  assign new_n787 = ~new_n687 & ~new_n782;
  assign new_n788 = ~new_n783 & ~new_n787;
  assign new_n789 = ~new_n687 & new_n788;
  assign new_n790 = ~new_n786 & ~new_n789;
  assign new_n791 = new_n786 & new_n789;
  assign new_n792 = ~new_n790 & ~new_n791;
  assign new_n793 = ~new_n690 & ~new_n792;
  assign new_n794 = ~new_n690 & new_n793;
  assign new_n795 = ~new_n776 & ~new_n794;
  assign new_n796 = new_n690 & ~new_n782;
  assign new_n797 = new_n690 & new_n796;
  assign new_n798 = new_n687 & ~new_n788;
  assign new_n799 = ~new_n789 & ~new_n798;
  assign new_n800 = ~new_n690 & ~new_n799;
  assign new_n801 = ~new_n690 & new_n800;
  assign new_n802 = ~new_n797 & ~new_n801;
  assign new_n803 = new_n695 & new_n802;
  assign new_n804 = ~new_n795 & ~new_n803;
  assign new_n805 = new_n795 & new_n803;
  assign new_n806 = ~new_n804 & ~new_n805;
  assign new_n807 = ~new_n675 & ~new_n806;
  assign new_n808 = ~new_n675 & new_n807;
  assign new_n809 = ~new_n774 & ~new_n808;
  assign new_n810 = \V223(1)  & ~new_n545;
  assign new_n811 = new_n567 & new_n810;
  assign new_n812 = \V183(1)  & new_n545;
  assign new_n813 = ~new_n567 & new_n812;
  assign new_n814 = ~new_n811 & ~new_n813;
  assign new_n815 = new_n704 & ~new_n814;
  assign new_n816 = new_n534 & new_n815;
  assign new_n817 = ~new_n542 & new_n816;
  assign new_n818 = ~new_n578 & new_n817;
  assign new_n819 = ~new_n662 & new_n818;
  assign new_n820 = new_n661 & new_n819;
  assign new_n821 = \V32(1)  & new_n662;
  assign new_n822 = ~new_n661 & new_n821;
  assign \V1213(1)  = new_n820 | new_n822;
  assign new_n824 = ~new_n809 & ~\V1213(1) ;
  assign new_n825 = new_n809 & \V1213(1) ;
  assign new_n826 = ~new_n824 & ~new_n825;
  assign new_n827 = new_n753 & new_n754;
  assign new_n828 = ~new_n752 & new_n753;
  assign new_n829 = ~new_n752 & new_n754;
  assign new_n830 = ~new_n827 & ~new_n828;
  assign new_n831 = ~new_n829 & new_n830;
  assign new_n832 = new_n754 & new_n831;
  assign new_n833 = ~new_n754 & ~new_n831;
  assign new_n834 = ~new_n832 & ~new_n833;
  assign new_n835 = new_n747 & ~new_n760;
  assign new_n836 = ~new_n746 & new_n747;
  assign new_n837 = ~new_n746 & ~new_n760;
  assign new_n838 = ~new_n835 & ~new_n836;
  assign new_n839 = ~new_n837 & new_n838;
  assign new_n840 = ~new_n834 & new_n839;
  assign new_n841 = new_n834 & ~new_n839;
  assign new_n842 = ~new_n840 & ~new_n841;
  assign new_n843 = new_n741 & ~new_n766;
  assign new_n844 = ~new_n740 & new_n741;
  assign new_n845 = ~new_n740 & ~new_n766;
  assign new_n846 = ~new_n843 & ~new_n844;
  assign new_n847 = ~new_n845 & new_n846;
  assign new_n848 = ~new_n842 & new_n847;
  assign new_n849 = new_n842 & ~new_n847;
  assign new_n850 = ~new_n848 & ~new_n849;
  assign new_n851 = new_n675 & ~new_n850;
  assign new_n852 = new_n675 & new_n851;
  assign new_n853 = new_n690 & ~new_n850;
  assign new_n854 = new_n690 & new_n853;
  assign new_n855 = ~new_n785 & ~new_n850;
  assign new_n856 = new_n785 & new_n850;
  assign new_n857 = ~new_n855 & ~new_n856;
  assign new_n858 = ~new_n791 & ~new_n857;
  assign new_n859 = new_n791 & new_n857;
  assign new_n860 = ~new_n858 & ~new_n859;
  assign new_n861 = ~new_n690 & ~new_n860;
  assign new_n862 = ~new_n690 & new_n861;
  assign new_n863 = ~new_n854 & ~new_n862;
  assign new_n864 = ~new_n805 & ~new_n863;
  assign new_n865 = new_n805 & new_n863;
  assign new_n866 = ~new_n864 & ~new_n865;
  assign new_n867 = ~new_n675 & ~new_n866;
  assign new_n868 = ~new_n675 & new_n867;
  assign new_n869 = ~new_n852 & ~new_n868;
  assign new_n870 = \V223(0)  & ~new_n545;
  assign new_n871 = new_n567 & new_n870;
  assign new_n872 = \V183(0)  & new_n545;
  assign new_n873 = ~new_n567 & new_n872;
  assign new_n874 = ~new_n871 & ~new_n873;
  assign new_n875 = new_n704 & ~new_n874;
  assign new_n876 = new_n534 & new_n875;
  assign new_n877 = ~new_n542 & new_n876;
  assign new_n878 = ~new_n578 & new_n877;
  assign new_n879 = ~new_n662 & new_n878;
  assign new_n880 = new_n661 & new_n879;
  assign new_n881 = \V32(0)  & new_n662;
  assign new_n882 = ~new_n661 & new_n881;
  assign \V1213(0)  = new_n880 | new_n882;
  assign new_n884 = ~new_n869 & ~\V1213(0) ;
  assign new_n885 = new_n869 & \V1213(0) ;
  assign new_n886 = ~new_n884 & ~new_n885;
  assign new_n887 = new_n675 & ~new_n782;
  assign new_n888 = new_n675 & new_n887;
  assign new_n889 = ~new_n695 & ~new_n802;
  assign new_n890 = ~new_n803 & ~new_n889;
  assign new_n891 = ~new_n675 & ~new_n890;
  assign new_n892 = ~new_n675 & new_n891;
  assign new_n893 = ~new_n888 & ~new_n892;
  assign new_n894 = \V223(2)  & ~new_n545;
  assign new_n895 = new_n567 & new_n894;
  assign new_n896 = \V183(2)  & new_n545;
  assign new_n897 = ~new_n567 & new_n896;
  assign new_n898 = ~new_n895 & ~new_n897;
  assign new_n899 = new_n704 & ~new_n898;
  assign new_n900 = new_n534 & new_n899;
  assign new_n901 = ~new_n542 & new_n900;
  assign new_n902 = ~new_n578 & new_n901;
  assign new_n903 = ~new_n662 & new_n902;
  assign new_n904 = new_n661 & new_n903;
  assign new_n905 = \V32(2)  & new_n662;
  assign new_n906 = ~new_n661 & new_n905;
  assign \V1213(2)  = new_n904 | new_n906;
  assign new_n908 = ~new_n893 & ~\V1213(2) ;
  assign new_n909 = new_n893 & \V1213(2) ;
  assign new_n910 = ~new_n908 & ~new_n909;
  assign new_n911 = ~\V288(0)  & ~\V288(1) ;
  assign new_n912 = ~new_n673 & new_n716;
  assign new_n913 = new_n826 & new_n912;
  assign new_n914 = new_n886 & new_n913;
  assign new_n915 = new_n910 & new_n914;
  assign new_n916 = ~new_n911 & new_n915;
  assign new_n917 = new_n676 & ~new_n684;
  assign new_n918 = new_n676 & new_n917;
  assign new_n919 = ~new_n684 & new_n717;
  assign new_n920 = new_n717 & new_n919;
  assign new_n921 = ~new_n684 & ~new_n717;
  assign new_n922 = ~new_n717 & new_n921;
  assign new_n923 = ~new_n920 & ~new_n922;
  assign new_n924 = ~new_n676 & new_n923;
  assign new_n925 = ~new_n676 & new_n924;
  assign new_n926 = ~new_n918 & ~new_n925;
  assign new_n927 = ~\V1213(3)  & ~new_n926;
  assign new_n928 = \V1213(3)  & new_n926;
  assign new_n929 = ~new_n927 & ~new_n928;
  assign new_n930 = new_n676 & ~new_n766;
  assign new_n931 = new_n676 & new_n930;
  assign new_n932 = new_n717 & ~new_n766;
  assign new_n933 = new_n717 & new_n932;
  assign new_n934 = new_n684 & new_n734;
  assign new_n935 = ~new_n766 & ~new_n934;
  assign new_n936 = new_n766 & new_n934;
  assign new_n937 = ~new_n935 & ~new_n936;
  assign new_n938 = ~new_n684 & ~new_n734;
  assign new_n939 = ~new_n934 & ~new_n938;
  assign new_n940 = ~new_n684 & new_n939;
  assign new_n941 = ~new_n937 & ~new_n940;
  assign new_n942 = new_n937 & new_n940;
  assign new_n943 = ~new_n941 & ~new_n942;
  assign new_n944 = ~new_n717 & ~new_n943;
  assign new_n945 = ~new_n717 & new_n944;
  assign new_n946 = ~new_n933 & ~new_n945;
  assign new_n947 = new_n717 & ~new_n734;
  assign new_n948 = new_n717 & new_n947;
  assign new_n949 = new_n684 & ~new_n939;
  assign new_n950 = ~new_n940 & ~new_n949;
  assign new_n951 = ~new_n717 & ~new_n950;
  assign new_n952 = ~new_n717 & new_n951;
  assign new_n953 = ~new_n948 & ~new_n952;
  assign new_n954 = new_n923 & new_n953;
  assign new_n955 = ~new_n946 & ~new_n954;
  assign new_n956 = new_n946 & new_n954;
  assign new_n957 = ~new_n955 & ~new_n956;
  assign new_n958 = ~new_n676 & ~new_n957;
  assign new_n959 = ~new_n676 & new_n958;
  assign new_n960 = ~new_n931 & ~new_n959;
  assign new_n961 = ~\V1213(1)  & ~new_n960;
  assign new_n962 = \V1213(1)  & new_n960;
  assign new_n963 = ~new_n961 & ~new_n962;
  assign new_n964 = new_n676 & ~new_n842;
  assign new_n965 = new_n676 & new_n964;
  assign new_n966 = new_n717 & ~new_n842;
  assign new_n967 = new_n717 & new_n966;
  assign new_n968 = ~new_n842 & ~new_n936;
  assign new_n969 = new_n842 & new_n936;
  assign new_n970 = ~new_n968 & ~new_n969;
  assign new_n971 = ~new_n942 & ~new_n970;
  assign new_n972 = new_n942 & new_n970;
  assign new_n973 = ~new_n971 & ~new_n972;
  assign new_n974 = ~new_n717 & ~new_n973;
  assign new_n975 = ~new_n717 & new_n974;
  assign new_n976 = ~new_n967 & ~new_n975;
  assign new_n977 = ~new_n956 & ~new_n976;
  assign new_n978 = new_n956 & new_n976;
  assign new_n979 = ~new_n977 & ~new_n978;
  assign new_n980 = ~new_n676 & ~new_n979;
  assign new_n981 = ~new_n676 & new_n980;
  assign new_n982 = ~new_n965 & ~new_n981;
  assign new_n983 = ~\V1213(0)  & ~new_n982;
  assign new_n984 = \V1213(0)  & new_n982;
  assign new_n985 = ~new_n983 & ~new_n984;
  assign new_n986 = new_n676 & ~new_n734;
  assign new_n987 = new_n676 & new_n986;
  assign new_n988 = ~new_n923 & ~new_n953;
  assign new_n989 = ~new_n954 & ~new_n988;
  assign new_n990 = ~new_n676 & ~new_n989;
  assign new_n991 = ~new_n676 & new_n990;
  assign new_n992 = ~new_n987 & ~new_n991;
  assign new_n993 = ~\V1213(2)  & ~new_n992;
  assign new_n994 = \V1213(2)  & new_n992;
  assign new_n995 = ~new_n993 & ~new_n994;
  assign new_n996 = ~\V288(2)  & ~\V288(3) ;
  assign new_n997 = ~new_n673 & new_n929;
  assign new_n998 = new_n963 & new_n997;
  assign new_n999 = new_n985 & new_n998;
  assign new_n1000 = new_n995 & new_n999;
  assign new_n1001 = ~new_n996 & new_n1000;
  assign new_n1002 = new_n677 & ~new_n681;
  assign new_n1003 = new_n677 & new_n1002;
  assign new_n1004 = ~new_n681 & new_n718;
  assign new_n1005 = new_n718 & new_n1004;
  assign new_n1006 = ~new_n681 & ~new_n718;
  assign new_n1007 = ~new_n718 & new_n1006;
  assign new_n1008 = ~new_n1005 & ~new_n1007;
  assign new_n1009 = ~new_n677 & new_n1008;
  assign new_n1010 = ~new_n677 & new_n1009;
  assign new_n1011 = ~new_n1003 & ~new_n1010;
  assign new_n1012 = ~\V1213(3)  & ~new_n1011;
  assign new_n1013 = \V1213(3)  & new_n1011;
  assign new_n1014 = ~new_n1012 & ~new_n1013;
  assign new_n1015 = new_n677 & ~new_n760;
  assign new_n1016 = new_n677 & new_n1015;
  assign new_n1017 = new_n718 & ~new_n760;
  assign new_n1018 = new_n718 & new_n1017;
  assign new_n1019 = new_n681 & new_n727;
  assign new_n1020 = ~new_n760 & ~new_n1019;
  assign new_n1021 = new_n760 & new_n1019;
  assign new_n1022 = ~new_n1020 & ~new_n1021;
  assign new_n1023 = ~new_n681 & ~new_n727;
  assign new_n1024 = ~new_n1019 & ~new_n1023;
  assign new_n1025 = ~new_n681 & new_n1024;
  assign new_n1026 = ~new_n1022 & ~new_n1025;
  assign new_n1027 = new_n1022 & new_n1025;
  assign new_n1028 = ~new_n1026 & ~new_n1027;
  assign new_n1029 = ~new_n718 & ~new_n1028;
  assign new_n1030 = ~new_n718 & new_n1029;
  assign new_n1031 = ~new_n1018 & ~new_n1030;
  assign new_n1032 = new_n718 & ~new_n727;
  assign new_n1033 = new_n718 & new_n1032;
  assign new_n1034 = new_n681 & ~new_n1024;
  assign new_n1035 = ~new_n1025 & ~new_n1034;
  assign new_n1036 = ~new_n718 & ~new_n1035;
  assign new_n1037 = ~new_n718 & new_n1036;
  assign new_n1038 = ~new_n1033 & ~new_n1037;
  assign new_n1039 = new_n1008 & new_n1038;
  assign new_n1040 = ~new_n1031 & ~new_n1039;
  assign new_n1041 = new_n1031 & new_n1039;
  assign new_n1042 = ~new_n1040 & ~new_n1041;
  assign new_n1043 = ~new_n677 & ~new_n1042;
  assign new_n1044 = ~new_n677 & new_n1043;
  assign new_n1045 = ~new_n1016 & ~new_n1044;
  assign new_n1046 = ~\V1213(1)  & ~new_n1045;
  assign new_n1047 = \V1213(1)  & new_n1045;
  assign new_n1048 = ~new_n1046 & ~new_n1047;
  assign new_n1049 = new_n677 & ~new_n834;
  assign new_n1050 = new_n677 & new_n1049;
  assign new_n1051 = new_n718 & ~new_n834;
  assign new_n1052 = new_n718 & new_n1051;
  assign new_n1053 = ~new_n834 & ~new_n1021;
  assign new_n1054 = new_n834 & new_n1021;
  assign new_n1055 = ~new_n1053 & ~new_n1054;
  assign new_n1056 = ~new_n1027 & ~new_n1055;
  assign new_n1057 = new_n1027 & new_n1055;
  assign new_n1058 = ~new_n1056 & ~new_n1057;
  assign new_n1059 = ~new_n718 & ~new_n1058;
  assign new_n1060 = ~new_n718 & new_n1059;
  assign new_n1061 = ~new_n1052 & ~new_n1060;
  assign new_n1062 = ~new_n1041 & ~new_n1061;
  assign new_n1063 = new_n1041 & new_n1061;
  assign new_n1064 = ~new_n1062 & ~new_n1063;
  assign new_n1065 = ~new_n677 & ~new_n1064;
  assign new_n1066 = ~new_n677 & new_n1065;
  assign new_n1067 = ~new_n1050 & ~new_n1066;
  assign new_n1068 = ~\V1213(0)  & ~new_n1067;
  assign new_n1069 = \V1213(0)  & new_n1067;
  assign new_n1070 = ~new_n1068 & ~new_n1069;
  assign new_n1071 = new_n677 & ~new_n727;
  assign new_n1072 = new_n677 & new_n1071;
  assign new_n1073 = ~new_n1008 & ~new_n1038;
  assign new_n1074 = ~new_n1039 & ~new_n1073;
  assign new_n1075 = ~new_n677 & ~new_n1074;
  assign new_n1076 = ~new_n677 & new_n1075;
  assign new_n1077 = ~new_n1072 & ~new_n1076;
  assign new_n1078 = ~\V1213(2)  & ~new_n1077;
  assign new_n1079 = \V1213(2)  & new_n1077;
  assign new_n1080 = ~new_n1078 & ~new_n1079;
  assign new_n1081 = ~\V288(4)  & ~\V288(5) ;
  assign new_n1082 = ~new_n673 & new_n1014;
  assign new_n1083 = new_n1048 & new_n1082;
  assign new_n1084 = new_n1070 & new_n1083;
  assign new_n1085 = new_n1080 & new_n1084;
  assign new_n1086 = ~new_n1081 & new_n1085;
  assign new_n1087 = ~new_n673 & ~\V1213(3) ;
  assign new_n1088 = ~\V1213(1)  & new_n1087;
  assign new_n1089 = ~\V1213(0)  & new_n1088;
  assign new_n1090 = ~\V1213(2)  & new_n1089;
  assign new_n1091 = ~new_n754 & new_n1090;
  assign new_n1092 = ~new_n673 & \V1213(2) ;
  assign new_n1093 = ~\V1213(1)  & new_n1092;
  assign new_n1094 = ~\V1213(0)  & new_n1093;
  assign new_n1095 = ~\V1213(3)  & new_n1094;
  assign new_n1096 = \V288(6)  & new_n1095;
  assign new_n1097 = \V288(7)  & new_n1096;
  assign new_n1098 = new_n681 & ~\V1213(3) ;
  assign new_n1099 = ~new_n681 & \V1213(3) ;
  assign new_n1100 = ~new_n1098 & ~new_n1099;
  assign new_n1101 = ~\V1213(1)  & ~new_n1022;
  assign new_n1102 = \V1213(1)  & new_n1022;
  assign new_n1103 = ~new_n1101 & ~new_n1102;
  assign new_n1104 = ~\V1213(0)  & ~new_n1055;
  assign new_n1105 = \V1213(0)  & new_n1055;
  assign new_n1106 = ~new_n1104 & ~new_n1105;
  assign new_n1107 = ~\V1213(2)  & ~new_n1024;
  assign new_n1108 = \V1213(2)  & new_n1024;
  assign new_n1109 = ~new_n1107 & ~new_n1108;
  assign new_n1110 = ~new_n673 & new_n1100;
  assign new_n1111 = new_n1103 & new_n1110;
  assign new_n1112 = new_n1106 & new_n1111;
  assign new_n1113 = new_n1109 & new_n1112;
  assign new_n1114 = new_n753 & new_n1113;
  assign new_n1115 = new_n684 & ~\V1213(3) ;
  assign new_n1116 = ~new_n684 & \V1213(3) ;
  assign new_n1117 = ~new_n1115 & ~new_n1116;
  assign new_n1118 = ~\V1213(1)  & ~new_n937;
  assign new_n1119 = \V1213(1)  & new_n937;
  assign new_n1120 = ~new_n1118 & ~new_n1119;
  assign new_n1121 = ~\V1213(0)  & ~new_n970;
  assign new_n1122 = \V1213(0)  & new_n970;
  assign new_n1123 = ~new_n1121 & ~new_n1122;
  assign new_n1124 = ~\V1213(2)  & ~new_n939;
  assign new_n1125 = \V1213(2)  & new_n939;
  assign new_n1126 = ~new_n1124 & ~new_n1125;
  assign new_n1127 = ~new_n673 & new_n1117;
  assign new_n1128 = new_n1120 & new_n1127;
  assign new_n1129 = new_n1123 & new_n1128;
  assign new_n1130 = new_n1126 & new_n1129;
  assign new_n1131 = new_n747 & new_n1130;
  assign new_n1132 = new_n687 & ~\V1213(3) ;
  assign new_n1133 = ~new_n687 & \V1213(3) ;
  assign new_n1134 = ~new_n1132 & ~new_n1133;
  assign new_n1135 = ~new_n786 & ~\V1213(1) ;
  assign new_n1136 = new_n786 & \V1213(1) ;
  assign new_n1137 = ~new_n1135 & ~new_n1136;
  assign new_n1138 = ~new_n857 & ~\V1213(0) ;
  assign new_n1139 = new_n857 & \V1213(0) ;
  assign new_n1140 = ~new_n1138 & ~new_n1139;
  assign new_n1141 = ~new_n788 & ~\V1213(2) ;
  assign new_n1142 = new_n788 & \V1213(2) ;
  assign new_n1143 = ~new_n1141 & ~new_n1142;
  assign new_n1144 = ~new_n673 & new_n1134;
  assign new_n1145 = new_n1137 & new_n1144;
  assign new_n1146 = new_n1140 & new_n1145;
  assign new_n1147 = new_n1143 & new_n1146;
  assign new_n1148 = new_n741 & new_n1147;
  assign new_n1149 = new_n674 & ~new_n916;
  assign new_n1150 = ~new_n1001 & new_n1149;
  assign new_n1151 = ~new_n1086 & new_n1150;
  assign new_n1152 = ~new_n1091 & new_n1151;
  assign new_n1153 = ~new_n1097 & new_n1152;
  assign new_n1154 = ~new_n1114 & new_n1153;
  assign new_n1155 = ~new_n1131 & new_n1154;
  assign V356 = ~new_n1148 & new_n1155;
  assign new_n1157 = ~new_n695 & ~\V1213(3) ;
  assign new_n1158 = new_n695 & \V1213(3) ;
  assign new_n1159 = ~new_n1157 & ~new_n1158;
  assign new_n1160 = ~new_n795 & ~\V1213(1) ;
  assign new_n1161 = new_n795 & \V1213(1) ;
  assign new_n1162 = ~new_n1160 & ~new_n1161;
  assign new_n1163 = ~new_n863 & ~\V1213(0) ;
  assign new_n1164 = new_n863 & \V1213(0) ;
  assign new_n1165 = ~new_n1163 & ~new_n1164;
  assign new_n1166 = ~new_n802 & ~\V1213(2) ;
  assign new_n1167 = new_n802 & \V1213(2) ;
  assign new_n1168 = ~new_n1166 & ~new_n1167;
  assign new_n1169 = ~new_n673 & new_n1159;
  assign new_n1170 = new_n1162 & new_n1169;
  assign new_n1171 = new_n1165 & new_n1170;
  assign new_n1172 = new_n1168 & new_n1171;
  assign new_n1173 = \V288(0)  & new_n1172;
  assign new_n1174 = ~\V1213(3)  & ~new_n923;
  assign new_n1175 = \V1213(3)  & new_n923;
  assign new_n1176 = ~new_n1174 & ~new_n1175;
  assign new_n1177 = ~\V1213(1)  & ~new_n946;
  assign new_n1178 = \V1213(1)  & new_n946;
  assign new_n1179 = ~new_n1177 & ~new_n1178;
  assign new_n1180 = ~\V1213(0)  & ~new_n976;
  assign new_n1181 = \V1213(0)  & new_n976;
  assign new_n1182 = ~new_n1180 & ~new_n1181;
  assign new_n1183 = ~\V1213(2)  & ~new_n953;
  assign new_n1184 = \V1213(2)  & new_n953;
  assign new_n1185 = ~new_n1183 & ~new_n1184;
  assign new_n1186 = ~new_n673 & new_n1176;
  assign new_n1187 = new_n1179 & new_n1186;
  assign new_n1188 = new_n1182 & new_n1187;
  assign new_n1189 = new_n1185 & new_n1188;
  assign new_n1190 = \V288(2)  & new_n1189;
  assign new_n1191 = ~\V1213(3)  & ~new_n1008;
  assign new_n1192 = \V1213(3)  & new_n1008;
  assign new_n1193 = ~new_n1191 & ~new_n1192;
  assign new_n1194 = ~\V1213(1)  & ~new_n1031;
  assign new_n1195 = \V1213(1)  & new_n1031;
  assign new_n1196 = ~new_n1194 & ~new_n1195;
  assign new_n1197 = ~\V1213(0)  & ~new_n1061;
  assign new_n1198 = \V1213(0)  & new_n1061;
  assign new_n1199 = ~new_n1197 & ~new_n1198;
  assign new_n1200 = ~\V1213(2)  & ~new_n1038;
  assign new_n1201 = \V1213(2)  & new_n1038;
  assign new_n1202 = ~new_n1200 & ~new_n1201;
  assign new_n1203 = ~new_n673 & new_n1193;
  assign new_n1204 = new_n1196 & new_n1203;
  assign new_n1205 = new_n1199 & new_n1204;
  assign new_n1206 = new_n1202 & new_n1205;
  assign new_n1207 = \V288(4)  & new_n1206;
  assign new_n1208 = ~new_n673 & \V1213(3) ;
  assign new_n1209 = ~\V1213(1)  & new_n1208;
  assign new_n1210 = ~\V1213(0)  & new_n1209;
  assign new_n1211 = ~\V1213(2)  & new_n1210;
  assign new_n1212 = \V288(6)  & new_n1211;
  assign new_n1213 = ~new_n673 & ~\V1213(1) ;
  assign new_n1214 = ~\V1213(0)  & new_n1213;
  assign new_n1215 = \V1213(2)  & new_n1214;
  assign new_n1216 = \V1213(3)  & new_n1215;
  assign new_n1217 = \V288(6)  & new_n1216;
  assign new_n1218 = \V288(7)  & new_n1217;
  assign new_n1219 = ~new_n681 & ~\V1213(3) ;
  assign new_n1220 = new_n681 & \V1213(3) ;
  assign new_n1221 = ~new_n1219 & ~new_n1220;
  assign new_n1222 = ~new_n760 & ~\V1213(1) ;
  assign new_n1223 = new_n760 & \V1213(1) ;
  assign new_n1224 = ~new_n1222 & ~new_n1223;
  assign new_n1225 = ~new_n834 & ~\V1213(0) ;
  assign new_n1226 = new_n834 & \V1213(0) ;
  assign new_n1227 = ~new_n1225 & ~new_n1226;
  assign new_n1228 = ~new_n727 & ~\V1213(2) ;
  assign new_n1229 = new_n727 & \V1213(2) ;
  assign new_n1230 = ~new_n1228 & ~new_n1229;
  assign new_n1231 = ~new_n673 & new_n1221;
  assign new_n1232 = new_n1224 & new_n1231;
  assign new_n1233 = new_n1227 & new_n1232;
  assign new_n1234 = new_n1230 & new_n1233;
  assign new_n1235 = new_n753 & new_n1234;
  assign new_n1236 = ~new_n684 & ~\V1213(3) ;
  assign new_n1237 = new_n684 & \V1213(3) ;
  assign new_n1238 = ~new_n1236 & ~new_n1237;
  assign new_n1239 = ~new_n766 & ~\V1213(1) ;
  assign new_n1240 = new_n766 & \V1213(1) ;
  assign new_n1241 = ~new_n1239 & ~new_n1240;
  assign new_n1242 = ~new_n842 & ~\V1213(0) ;
  assign new_n1243 = new_n842 & \V1213(0) ;
  assign new_n1244 = ~new_n1242 & ~new_n1243;
  assign new_n1245 = ~new_n734 & ~\V1213(2) ;
  assign new_n1246 = new_n734 & \V1213(2) ;
  assign new_n1247 = ~new_n1245 & ~new_n1246;
  assign new_n1248 = ~new_n673 & new_n1238;
  assign new_n1249 = new_n1241 & new_n1248;
  assign new_n1250 = new_n1244 & new_n1249;
  assign new_n1251 = new_n1247 & new_n1250;
  assign new_n1252 = new_n747 & new_n1251;
  assign new_n1253 = ~new_n687 & ~\V1213(3) ;
  assign new_n1254 = new_n687 & \V1213(3) ;
  assign new_n1255 = ~new_n1253 & ~new_n1254;
  assign new_n1256 = ~new_n772 & ~\V1213(1) ;
  assign new_n1257 = new_n772 & \V1213(1) ;
  assign new_n1258 = ~new_n1256 & ~new_n1257;
  assign new_n1259 = ~new_n850 & ~\V1213(0) ;
  assign new_n1260 = new_n850 & \V1213(0) ;
  assign new_n1261 = ~new_n1259 & ~new_n1260;
  assign new_n1262 = ~new_n782 & ~\V1213(2) ;
  assign new_n1263 = new_n782 & \V1213(2) ;
  assign new_n1264 = ~new_n1262 & ~new_n1263;
  assign new_n1265 = ~new_n673 & new_n1255;
  assign new_n1266 = new_n1258 & new_n1265;
  assign new_n1267 = new_n1261 & new_n1266;
  assign new_n1268 = new_n1264 & new_n1267;
  assign new_n1269 = new_n741 & new_n1268;
  assign new_n1270 = new_n534 & ~new_n1173;
  assign new_n1271 = ~new_n1190 & new_n1270;
  assign new_n1272 = ~new_n1207 & new_n1271;
  assign new_n1273 = ~new_n1212 & new_n1272;
  assign new_n1274 = ~new_n1218 & new_n1273;
  assign new_n1275 = ~new_n1235 & new_n1274;
  assign new_n1276 = ~new_n1252 & new_n1275;
  assign V357 = ~new_n1269 & new_n1276;
  assign V373 = \V10(0)  & \V13(0) ;
  assign new_n1279 = \V202(0)  & \V71(0) ;
  assign new_n1280 = ~\V13(0)  & new_n1279;
  assign new_n1281 = \V9(0)  & ~new_n1280;
  assign V789 = \V4(0)  & new_n1281;
  assign V1263 = \V9(0)  & \V4(0) ;
  assign V1259 = \V9(0)  & \V3(0) ;
  assign V1387 = \V9(0)  & \V8(0) ;
  assign V780 = \V9(0)  & \V6(0) ;
  assign V778 = \V9(0)  & \V5(0) ;
  assign V787 = \V7(0)  & \V9(0) ;
  assign new_n1289 = ~\V13(0)  & \V109(0) ;
  assign V1423 = \V1(0)  & \V9(0) ;
  assign V1431 = ~new_n1289 & V1423;
  assign V1258 = \V9(0)  & \V2(0) ;
  assign new_n1293 = ~V787 & ~V1431;
  assign new_n1294 = ~V1258 & new_n1293;
  assign new_n1295 = ~V1423 & new_n1294;
  assign new_n1296 = ~V1387 & ~V780;
  assign new_n1297 = ~V778 & new_n1296;
  assign new_n1298 = ~V789 & ~V1263;
  assign new_n1299 = ~V1259 & new_n1298;
  assign new_n1300 = new_n1297 & new_n1299;
  assign \V375(0)  = ~new_n1295 | ~new_n1300;
  assign new_n1302 = \V203(0)  & \V165(1) ;
  assign new_n1303 = ~\V165(0)  & new_n1302;
  assign new_n1304 = \V165(2)  & new_n1303;
  assign new_n1305 = ~\V35(0)  & ~new_n1304;
  assign V377 = \V203(0)  & ~new_n1305;
  assign new_n1307 = \V243(0)  & \V244(0) ;
  assign new_n1308 = \V245(0)  & new_n1307;
  assign new_n1309 = \V246(0)  & new_n1308;
  assign new_n1310 = \V165(0)  & ~\V165(2) ;
  assign new_n1311 = \V165(1)  & new_n1310;
  assign new_n1312 = \V240(0)  & ~new_n1311;
  assign V1719 = ~\V172(0)  & new_n1312;
  assign new_n1314 = ~\V248(0)  & new_n1309;
  assign new_n1315 = V1719 & new_n1314;
  assign new_n1316 = \V247(0)  & new_n1315;
  assign new_n1317 = new_n534 & ~new_n1091;
  assign new_n1318 = ~new_n1212 & new_n1317;
  assign new_n1319 = new_n534 & ~new_n1097;
  assign new_n1320 = ~new_n1218 & new_n1319;
  assign new_n1321 = new_n1318 & new_n1320;
  assign new_n1322 = \V288(6)  & ~new_n1321;
  assign new_n1323 = \V288(7)  & new_n1322;
  assign new_n1324 = new_n534 & ~new_n1001;
  assign new_n1325 = ~new_n1190 & new_n1324;
  assign new_n1326 = new_n534 & ~new_n1131;
  assign new_n1327 = ~new_n1252 & new_n1326;
  assign new_n1328 = new_n1325 & new_n1327;
  assign new_n1329 = new_n747 & ~new_n1328;
  assign new_n1330 = new_n534 & ~new_n916;
  assign new_n1331 = ~new_n1173 & new_n1330;
  assign new_n1332 = new_n534 & ~new_n1148;
  assign new_n1333 = ~new_n1269 & new_n1332;
  assign new_n1334 = new_n1331 & new_n1333;
  assign new_n1335 = new_n741 & ~new_n1334;
  assign new_n1336 = new_n534 & ~new_n1086;
  assign new_n1337 = ~new_n1207 & new_n1336;
  assign new_n1338 = new_n534 & ~new_n1114;
  assign new_n1339 = ~new_n1235 & new_n1338;
  assign new_n1340 = new_n1337 & new_n1339;
  assign new_n1341 = new_n753 & ~new_n1340;
  assign new_n1342 = ~new_n1335 & ~new_n1341;
  assign new_n1343 = ~new_n1323 & ~new_n1329;
  assign new_n1344 = new_n1342 & new_n1343;
  assign new_n1345 = \V239(3)  & ~new_n545;
  assign new_n1346 = new_n567 & new_n1345;
  assign new_n1347 = \V199(3)  & new_n545;
  assign new_n1348 = ~new_n567 & new_n1347;
  assign new_n1349 = ~new_n1346 & ~new_n1348;
  assign new_n1350 = ~new_n557 & ~new_n1349;
  assign new_n1351 = new_n534 & new_n1350;
  assign new_n1352 = ~new_n542 & new_n1351;
  assign new_n1353 = ~new_n578 & new_n1352;
  assign new_n1354 = ~new_n578 & new_n1353;
  assign new_n1355 = \V32(10)  & new_n583;
  assign new_n1356 = new_n578 & new_n1355;
  assign new_n1357 = new_n578 & new_n1356;
  assign new_n1358 = ~new_n1354 & ~new_n1357;
  assign new_n1359 = ~new_n662 & ~new_n1358;
  assign new_n1360 = new_n661 & new_n1359;
  assign new_n1361 = \V88(0)  & new_n662;
  assign new_n1362 = ~new_n661 & new_n1361;
  assign \V1243(8)  = new_n1360 | new_n1362;
  assign new_n1364 = \V239(2)  & ~new_n545;
  assign new_n1365 = new_n567 & new_n1364;
  assign new_n1366 = \V199(2)  & new_n545;
  assign new_n1367 = ~new_n567 & new_n1366;
  assign new_n1368 = ~new_n1365 & ~new_n1367;
  assign new_n1369 = ~new_n557 & ~new_n1368;
  assign new_n1370 = new_n534 & new_n1369;
  assign new_n1371 = ~new_n542 & new_n1370;
  assign new_n1372 = ~new_n578 & new_n1371;
  assign new_n1373 = ~new_n578 & new_n1372;
  assign new_n1374 = \V32(9)  & new_n583;
  assign new_n1375 = new_n578 & new_n1374;
  assign new_n1376 = new_n578 & new_n1375;
  assign new_n1377 = ~new_n1373 & ~new_n1376;
  assign new_n1378 = ~new_n662 & ~new_n1377;
  assign new_n1379 = new_n661 & new_n1378;
  assign new_n1380 = \V84(5)  & new_n662;
  assign new_n1381 = ~new_n661 & new_n1380;
  assign \V1243(7)  = new_n1379 | new_n1381;
  assign new_n1383 = \V239(4)  & ~new_n545;
  assign new_n1384 = new_n567 & new_n1383;
  assign new_n1385 = \V199(4)  & new_n545;
  assign new_n1386 = ~new_n567 & new_n1385;
  assign new_n1387 = ~new_n1384 & ~new_n1386;
  assign new_n1388 = ~new_n557 & ~new_n1387;
  assign new_n1389 = new_n534 & new_n1388;
  assign new_n1390 = ~new_n542 & new_n1389;
  assign new_n1391 = ~new_n578 & new_n1390;
  assign new_n1392 = ~new_n578 & new_n1391;
  assign new_n1393 = \V32(11)  & new_n583;
  assign new_n1394 = new_n578 & new_n1393;
  assign new_n1395 = new_n578 & new_n1394;
  assign new_n1396 = ~new_n1392 & ~new_n1395;
  assign new_n1397 = ~new_n662 & ~new_n1396;
  assign new_n1398 = new_n661 & new_n1397;
  assign new_n1399 = \V88(1)  & new_n662;
  assign new_n1400 = ~new_n661 & new_n1399;
  assign \V1243(9)  = new_n1398 | new_n1400;
  assign new_n1402 = ~\V248(0)  & ~new_n1344;
  assign new_n1403 = \V1243(8)  & new_n1402;
  assign new_n1404 = \V1243(7)  & new_n1403;
  assign new_n1405 = \V1243(9)  & new_n1404;
  assign new_n1406 = V1719 & new_n1405;
  assign new_n1407 = \V199(4)  & \V199(2) ;
  assign new_n1408 = \V199(0)  & new_n1407;
  assign new_n1409 = \V194(3)  & new_n1408;
  assign new_n1410 = \V194(1)  & new_n1409;
  assign new_n1411 = \V194(2)  & new_n1410;
  assign new_n1412 = \V194(4)  & new_n1411;
  assign new_n1413 = \V199(1)  & new_n1412;
  assign new_n1414 = \V199(3)  & new_n1413;
  assign new_n1415 = ~\V248(0)  & new_n1414;
  assign new_n1416 = V1719 & new_n1415;
  assign new_n1417 = ~new_n1316 & ~new_n1406;
  assign \V393(0)  = new_n1416 | ~new_n1417;
  assign new_n1419 = ~V763 & ~new_n627;
  assign new_n1420 = \V802(0)  & ~new_n1419;
  assign new_n1421 = ~new_n540 & ~new_n567;
  assign new_n1422 = \V802(0)  & new_n1421;
  assign new_n1423 = \V66(0)  & ~new_n1311;
  assign new_n1424 = V763 & new_n1423;
  assign new_n1425 = ~\V215(0)  & new_n1424;
  assign new_n1426 = \V149(4)  & new_n644;
  assign new_n1427 = \V88(3)  & new_n603;
  assign new_n1428 = ~\V88(3)  & new_n616;
  assign new_n1429 = ~new_n1427 & ~new_n1428;
  assign new_n1430 = ~new_n627 & ~new_n1429;
  assign new_n1431 = ~new_n1426 & ~new_n1430;
  assign new_n1432 = ~\V174(0)  & ~new_n631;
  assign new_n1433 = ~new_n628 & new_n1431;
  assign new_n1434 = new_n1432 & new_n1433;
  assign new_n1435 = \V56(0)  & ~new_n1434;
  assign new_n1436 = new_n534 & new_n647;
  assign new_n1437 = ~new_n630 & new_n1436;
  assign new_n1438 = new_n648 & new_n1437;
  assign new_n1439 = \V802(0)  & ~new_n1438;
  assign new_n1440 = new_n627 & ~new_n1429;
  assign new_n1441 = ~new_n626 & ~new_n627;
  assign new_n1442 = new_n647 & ~new_n1440;
  assign new_n1443 = ~new_n1441 & new_n1442;
  assign new_n1444 = new_n534 & new_n1443;
  assign new_n1445 = \V59(0)  & ~new_n1444;
  assign new_n1446 = \V62(0)  & new_n628;
  assign new_n1447 = \V70(0)  & ~new_n534;
  assign new_n1448 = ~new_n1425 & ~new_n1435;
  assign new_n1449 = ~V1719 & ~new_n1422;
  assign new_n1450 = new_n1448 & new_n1449;
  assign new_n1451 = ~new_n1446 & ~new_n1447;
  assign new_n1452 = ~new_n1439 & ~new_n1445;
  assign new_n1453 = new_n1451 & new_n1452;
  assign \V423(0)  = ~new_n1450 | ~new_n1453;
  assign new_n1455 = \V248(0)  & V1719;
  assign new_n1456 = ~\V423(0)  & ~new_n1455;
  assign new_n1457 = ~\V165(7)  & new_n1311;
  assign new_n1458 = V1719 & new_n1457;
  assign new_n1459 = \V302(0)  & V1719;
  assign new_n1460 = new_n1304 & V1719;
  assign new_n1461 = ~\V214(0)  & ~new_n1420;
  assign new_n1462 = ~new_n1456 & new_n1461;
  assign new_n1463 = ~\V43(0)  & new_n1462;
  assign new_n1464 = ~new_n1458 & new_n1463;
  assign new_n1465 = ~new_n1459 & new_n1464;
  assign new_n1466 = ~new_n1416 & new_n1465;
  assign new_n1467 = ~new_n1406 & new_n1466;
  assign new_n1468 = ~new_n1460 & new_n1467;
  assign \V398(0)  = new_n1316 | ~new_n1468;
  assign new_n1470 = \V56(0)  & ~new_n1431;
  assign new_n1471 = \V59(0)  & ~new_n1443;
  assign new_n1472 = ~new_n1446 & ~new_n1470;
  assign new_n1473 = ~new_n1471 & new_n1472;
  assign new_n1474 = ~\V16(0)  & \V15(0) ;
  assign new_n1475 = \V16(0)  & \V15(0) ;
  assign \V1757(0)  = new_n1474 | new_n1475;
  assign new_n1477 = ~new_n1311 & ~new_n1473;
  assign \V410(0)  = \V1757(0)  | ~new_n1477;
  assign new_n1479 = \V215(0)  & \V66(0) ;
  assign new_n1480 = ~\V32(2)  & ~new_n782;
  assign new_n1481 = \V32(2)  & new_n782;
  assign new_n1482 = ~new_n1480 & ~new_n1481;
  assign new_n1483 = ~\V32(0)  & ~new_n850;
  assign new_n1484 = \V32(0)  & new_n850;
  assign new_n1485 = ~new_n1483 & ~new_n1484;
  assign new_n1486 = ~\V32(1)  & ~new_n772;
  assign new_n1487 = \V32(1)  & new_n772;
  assign new_n1488 = ~new_n1486 & ~new_n1487;
  assign new_n1489 = new_n1482 & new_n1485;
  assign new_n1490 = \V32(3)  & new_n1489;
  assign new_n1491 = new_n687 & new_n1490;
  assign new_n1492 = new_n1488 & new_n1491;
  assign new_n1493 = \V32(1)  & new_n1485;
  assign new_n1494 = new_n772 & new_n1493;
  assign new_n1495 = new_n782 & new_n1488;
  assign new_n1496 = \V32(2)  & new_n1495;
  assign new_n1497 = new_n1485 & new_n1496;
  assign new_n1498 = ~new_n1484 & ~new_n1497;
  assign new_n1499 = ~new_n1492 & ~new_n1494;
  assign new_n1500 = new_n1498 & new_n1499;
  assign new_n1501 = \V66(0)  & V763;
  assign new_n1502 = ~\V149(4)  & new_n596;
  assign new_n1503 = \V149(6)  & new_n1502;
  assign new_n1504 = \V66(0)  & new_n1503;
  assign new_n1505 = ~new_n538 & ~new_n599;
  assign new_n1506 = \V802(0)  & ~new_n1505;
  assign new_n1507 = ~V763 & new_n1506;
  assign new_n1508 = \V802(0)  & new_n544;
  assign new_n1509 = ~\V174(0)  & new_n494;
  assign new_n1510 = ~\V149(4)  & new_n497;
  assign new_n1511 = \V149(6)  & new_n1510;
  assign new_n1512 = ~\V149(4)  & new_n492;
  assign new_n1513 = \V149(6)  & new_n1512;
  assign new_n1514 = ~\V149(6)  & new_n1512;
  assign new_n1515 = ~new_n1513 & ~new_n1514;
  assign new_n1516 = ~new_n1509 & ~new_n1511;
  assign new_n1517 = new_n1515 & new_n1516;
  assign new_n1518 = \V56(0)  & ~new_n1517;
  assign new_n1519 = ~new_n1508 & ~new_n1518;
  assign new_n1520 = ~new_n1501 & ~new_n1504;
  assign new_n1521 = ~new_n1507 & new_n1520;
  assign new_n1522 = new_n1519 & new_n1521;
  assign new_n1523 = ~new_n1500 & ~new_n1522;
  assign new_n1524 = ~\V88(2)  & \V88(3) ;
  assign new_n1525 = \V88(2)  & ~\V88(3) ;
  assign new_n1526 = ~new_n1524 & ~new_n1525;
  assign new_n1527 = \V88(1)  & ~\V88(0) ;
  assign new_n1528 = ~\V88(1)  & \V88(0) ;
  assign new_n1529 = ~new_n1527 & ~new_n1528;
  assign new_n1530 = ~new_n1526 & new_n1529;
  assign new_n1531 = new_n1526 & ~new_n1529;
  assign new_n1532 = ~new_n1530 & ~new_n1531;
  assign new_n1533 = \V84(5)  & ~\V84(4) ;
  assign new_n1534 = ~\V84(5)  & \V84(4) ;
  assign new_n1535 = ~new_n1533 & ~new_n1534;
  assign new_n1536 = \V84(3)  & ~\V84(2) ;
  assign new_n1537 = ~\V84(3)  & \V84(2) ;
  assign new_n1538 = ~new_n1536 & ~new_n1537;
  assign new_n1539 = ~new_n1535 & new_n1538;
  assign new_n1540 = new_n1535 & ~new_n1538;
  assign new_n1541 = ~new_n1539 & ~new_n1540;
  assign new_n1542 = ~new_n1532 & new_n1541;
  assign new_n1543 = new_n1532 & ~new_n1541;
  assign new_n1544 = ~new_n1542 & ~new_n1543;
  assign new_n1545 = \V94(1)  & new_n1544;
  assign new_n1546 = ~\V94(1)  & ~new_n1544;
  assign new_n1547 = ~new_n1545 & ~new_n1546;
  assign new_n1548 = \V84(1)  & ~\V84(0) ;
  assign new_n1549 = ~\V84(1)  & \V84(0) ;
  assign new_n1550 = ~new_n1548 & ~new_n1549;
  assign new_n1551 = \V78(5)  & ~\V78(4) ;
  assign new_n1552 = ~\V78(5)  & \V78(4) ;
  assign new_n1553 = ~new_n1551 & ~new_n1552;
  assign new_n1554 = ~new_n1550 & new_n1553;
  assign new_n1555 = new_n1550 & ~new_n1553;
  assign new_n1556 = ~new_n1554 & ~new_n1555;
  assign new_n1557 = ~\V78(2)  & \V78(3) ;
  assign new_n1558 = \V78(2)  & ~\V78(3) ;
  assign new_n1559 = ~new_n1557 & ~new_n1558;
  assign new_n1560 = \V78(1)  & ~\V78(0) ;
  assign new_n1561 = ~\V78(1)  & \V78(0) ;
  assign new_n1562 = ~new_n1560 & ~new_n1561;
  assign new_n1563 = ~new_n1559 & new_n1562;
  assign new_n1564 = new_n1559 & ~new_n1562;
  assign new_n1565 = ~new_n1563 & ~new_n1564;
  assign new_n1566 = ~new_n1556 & new_n1565;
  assign new_n1567 = new_n1556 & ~new_n1565;
  assign new_n1568 = ~new_n1566 & ~new_n1567;
  assign new_n1569 = \V94(0)  & new_n1568;
  assign new_n1570 = ~\V94(0)  & ~new_n1568;
  assign new_n1571 = ~new_n1569 & ~new_n1570;
  assign new_n1572 = ~new_n1547 & ~new_n1571;
  assign new_n1573 = ~\V149(3)  & new_n668;
  assign new_n1574 = new_n489 & new_n1573;
  assign new_n1575 = \V149(4)  & new_n1574;
  assign new_n1576 = \V149(6)  & new_n1575;
  assign new_n1577 = ~new_n598 & ~new_n1514;
  assign new_n1578 = ~new_n1576 & new_n1577;
  assign new_n1579 = \V56(0)  & ~new_n1578;
  assign new_n1580 = ~new_n544 & ~new_n599;
  assign new_n1581 = ~new_n538 & new_n1580;
  assign new_n1582 = \V802(0)  & ~new_n1581;
  assign new_n1583 = ~new_n1579 & ~new_n1582;
  assign new_n1584 = ~new_n1572 & ~new_n1583;
  assign new_n1585 = \V56(0)  & \V172(0) ;
  assign new_n1586 = \V207(0)  & ~new_n1585;
  assign new_n1587 = ~\V43(0)  & ~\V214(0) ;
  assign new_n1588 = new_n534 & new_n1587;
  assign new_n1589 = ~new_n1479 & new_n1588;
  assign new_n1590 = ~new_n1523 & new_n1589;
  assign new_n1591 = ~\V1757(0)  & new_n1590;
  assign new_n1592 = ~new_n1420 & new_n1591;
  assign new_n1593 = ~new_n1584 & new_n1592;
  assign new_n1594 = ~new_n1586 & new_n1593;
  assign new_n1595 = \V423(0)  & new_n1594;
  assign new_n1596 = ~new_n1458 & new_n1595;
  assign new_n1597 = ~new_n1459 & new_n1596;
  assign new_n1598 = ~new_n1416 & new_n1597;
  assign new_n1599 = ~new_n1406 & new_n1598;
  assign new_n1600 = ~new_n1460 & new_n1599;
  assign V432 = ~new_n1316 & new_n1600;
  assign new_n1602 = \V56(0)  & new_n598;
  assign new_n1603 = \V241(0)  & ~new_n566;
  assign new_n1604 = ~new_n549 & ~new_n1603;
  assign new_n1605 = \V59(0)  & new_n540;
  assign new_n1606 = ~new_n1604 & new_n1605;
  assign new_n1607 = ~new_n538 & ~new_n549;
  assign new_n1608 = ~new_n537 & new_n1607;
  assign new_n1609 = new_n540 & ~new_n1608;
  assign new_n1610 = \V802(0)  & new_n1609;
  assign new_n1611 = ~\V270(0)  & ~new_n1610;
  assign new_n1612 = ~new_n1602 & ~new_n1606;
  assign new_n1613 = new_n1611 & new_n1612;
  assign new_n1614 = \V62(0)  & new_n598;
  assign new_n1615 = ~\V302(0)  & ~new_n1613;
  assign V630 = ~new_n1614 & new_n1615;
  assign \V435(0)  = V432 | V630;
  assign \V500(0)  = \V271(0)  | ~\V14(0) ;
  assign new_n1619 = \V59(0)  & new_n631;
  assign new_n1620 = new_n1514 & ~new_n1584;
  assign new_n1621 = ~new_n627 & new_n630;
  assign new_n1622 = ~new_n537 & ~new_n591;
  assign new_n1623 = ~new_n538 & ~new_n1620;
  assign new_n1624 = ~new_n1621 & new_n1623;
  assign new_n1625 = new_n1622 & new_n1624;
  assign new_n1626 = \V56(0)  & ~new_n1625;
  assign new_n1627 = \V62(0)  & new_n1513;
  assign new_n1628 = ~new_n1511 & ~new_n1513;
  assign new_n1629 = \V56(0)  & ~new_n1628;
  assign new_n1630 = ~new_n1627 & ~new_n1629;
  assign new_n1631 = ~new_n1619 & ~new_n1626;
  assign \V508(0)  = ~new_n1630 | ~new_n1631;
  assign new_n1633 = ~\V43(0)  & \V45(0) ;
  assign \V511(0)  = \V40(0)  | new_n1633;
  assign new_n1635 = \V42(0)  & ~\V44(0) ;
  assign new_n1636 = ~\V42(0)  & \V44(0) ;
  assign new_n1637 = ~new_n1635 & ~new_n1636;
  assign new_n1638 = \V39(0)  & ~\V38(0) ;
  assign new_n1639 = ~\V39(0)  & \V38(0) ;
  assign new_n1640 = ~new_n1638 & ~new_n1639;
  assign V512 = new_n1637 & new_n1640;
  assign new_n1642 = \V59(0)  & ~new_n627;
  assign new_n1643 = ~new_n626 & new_n1642;
  assign new_n1644 = \V56(0)  & new_n1426;
  assign new_n1645 = \V56(0)  & new_n1430;
  assign new_n1646 = \V59(0)  & new_n1440;
  assign new_n1647 = \V59(0)  & ~new_n647;
  assign new_n1648 = ~new_n1446 & ~new_n1643;
  assign new_n1649 = ~new_n1644 & new_n1648;
  assign new_n1650 = ~new_n1645 & new_n1649;
  assign new_n1651 = ~new_n1646 & new_n1650;
  assign new_n1652 = ~new_n1647 & new_n1651;
  assign new_n1653 = ~\V214(0)  & ~new_n1586;
  assign new_n1654 = ~new_n1652 & new_n1653;
  assign new_n1655 = ~new_n1311 & new_n1654;
  assign V527 = ~\V43(0)  & new_n1655;
  assign V537 = new_n538 & \V1213(0) ;
  assign V538 = new_n538 & \V1213(1) ;
  assign V539 = new_n538 & \V1213(2) ;
  assign V540 = new_n538 & \V1213(3) ;
  assign new_n1661 = \V257(6)  & ~new_n534;
  assign new_n1662 = ~new_n542 & new_n1661;
  assign new_n1663 = new_n557 & new_n1662;
  assign new_n1664 = \V223(4)  & ~new_n545;
  assign new_n1665 = new_n567 & new_n1664;
  assign new_n1666 = \V183(4)  & new_n545;
  assign new_n1667 = ~new_n567 & new_n1666;
  assign new_n1668 = ~new_n1665 & ~new_n1667;
  assign new_n1669 = new_n534 & ~new_n1668;
  assign new_n1670 = ~new_n542 & new_n1669;
  assign new_n1671 = ~new_n557 & new_n1670;
  assign new_n1672 = ~new_n1663 & ~new_n1671;
  assign new_n1673 = ~new_n578 & ~new_n1672;
  assign new_n1674 = ~new_n578 & new_n1673;
  assign new_n1675 = ~new_n662 & new_n1674;
  assign new_n1676 = new_n661 & new_n1675;
  assign new_n1677 = \V32(4)  & new_n662;
  assign new_n1678 = ~new_n661 & new_n1677;
  assign \V1213(4)  = new_n1676 | new_n1678;
  assign V541 = new_n538 & \V1213(4) ;
  assign new_n1681 = \V257(0)  & ~new_n534;
  assign new_n1682 = ~new_n542 & new_n1681;
  assign new_n1683 = new_n557 & new_n1682;
  assign new_n1684 = \V223(5)  & ~new_n545;
  assign new_n1685 = new_n567 & new_n1684;
  assign new_n1686 = \V183(5)  & new_n545;
  assign new_n1687 = ~new_n567 & new_n1686;
  assign new_n1688 = ~new_n1685 & ~new_n1687;
  assign new_n1689 = new_n534 & ~new_n1688;
  assign new_n1690 = ~new_n542 & new_n1689;
  assign new_n1691 = ~new_n557 & new_n1690;
  assign new_n1692 = ~new_n1683 & ~new_n1691;
  assign new_n1693 = ~new_n578 & ~new_n1692;
  assign new_n1694 = ~new_n578 & new_n1693;
  assign new_n1695 = new_n578 & ~new_n583;
  assign new_n1696 = new_n578 & new_n1695;
  assign new_n1697 = ~new_n1694 & ~new_n1696;
  assign new_n1698 = ~new_n662 & ~new_n1697;
  assign new_n1699 = new_n661 & new_n1698;
  assign new_n1700 = \V32(5)  & new_n662;
  assign new_n1701 = ~new_n661 & new_n1700;
  assign \V1213(5)  = new_n1699 | new_n1701;
  assign V542 = new_n538 & \V1213(5) ;
  assign new_n1704 = \V257(1)  & ~new_n534;
  assign new_n1705 = ~new_n542 & new_n1704;
  assign new_n1706 = new_n557 & new_n1705;
  assign new_n1707 = \V229(0)  & ~new_n545;
  assign new_n1708 = new_n567 & new_n1707;
  assign new_n1709 = \V189(0)  & new_n545;
  assign new_n1710 = ~new_n567 & new_n1709;
  assign new_n1711 = ~new_n1708 & ~new_n1710;
  assign new_n1712 = new_n534 & ~new_n1711;
  assign new_n1713 = ~new_n542 & new_n1712;
  assign new_n1714 = ~new_n557 & new_n1713;
  assign new_n1715 = ~new_n1706 & ~new_n1714;
  assign new_n1716 = ~new_n578 & ~new_n1715;
  assign new_n1717 = ~new_n578 & new_n1716;
  assign new_n1718 = new_n578 & new_n583;
  assign new_n1719 = new_n578 & new_n1718;
  assign new_n1720 = ~new_n1717 & ~new_n1719;
  assign new_n1721 = ~new_n662 & ~new_n1720;
  assign new_n1722 = new_n661 & new_n1721;
  assign new_n1723 = \V32(6)  & new_n662;
  assign new_n1724 = ~new_n661 & new_n1723;
  assign \V1213(6)  = new_n1722 | new_n1724;
  assign V543 = new_n538 & \V1213(6) ;
  assign new_n1727 = \V257(2)  & ~new_n534;
  assign new_n1728 = ~new_n542 & new_n1727;
  assign new_n1729 = new_n557 & new_n1728;
  assign new_n1730 = \V229(1)  & ~new_n545;
  assign new_n1731 = new_n567 & new_n1730;
  assign new_n1732 = \V189(1)  & new_n545;
  assign new_n1733 = ~new_n567 & new_n1732;
  assign new_n1734 = ~new_n1731 & ~new_n1733;
  assign new_n1735 = new_n534 & ~new_n1734;
  assign new_n1736 = ~new_n542 & new_n1735;
  assign new_n1737 = ~new_n557 & new_n1736;
  assign new_n1738 = ~new_n1729 & ~new_n1737;
  assign new_n1739 = ~new_n578 & ~new_n1738;
  assign new_n1740 = ~new_n578 & new_n1739;
  assign new_n1741 = \V32(0)  & ~new_n583;
  assign new_n1742 = ~new_n583 & new_n1741;
  assign new_n1743 = ~new_n583 & ~new_n1742;
  assign new_n1744 = new_n578 & ~new_n1743;
  assign new_n1745 = new_n578 & new_n1744;
  assign new_n1746 = ~new_n1740 & ~new_n1745;
  assign new_n1747 = ~new_n662 & ~new_n1746;
  assign new_n1748 = new_n661 & new_n1747;
  assign new_n1749 = \V32(7)  & new_n662;
  assign new_n1750 = ~new_n661 & new_n1749;
  assign \V1213(7)  = new_n1748 | new_n1750;
  assign V544 = new_n538 & \V1213(7) ;
  assign new_n1753 = \V257(3)  & ~new_n534;
  assign new_n1754 = ~new_n542 & new_n1753;
  assign new_n1755 = new_n557 & new_n1754;
  assign new_n1756 = \V229(2)  & ~new_n545;
  assign new_n1757 = new_n567 & new_n1756;
  assign new_n1758 = \V189(2)  & new_n545;
  assign new_n1759 = ~new_n567 & new_n1758;
  assign new_n1760 = ~new_n1757 & ~new_n1759;
  assign new_n1761 = new_n534 & ~new_n1760;
  assign new_n1762 = ~new_n542 & new_n1761;
  assign new_n1763 = ~new_n557 & new_n1762;
  assign new_n1764 = ~new_n1755 & ~new_n1763;
  assign new_n1765 = ~new_n578 & ~new_n1764;
  assign new_n1766 = ~new_n578 & new_n1765;
  assign new_n1767 = \V32(1)  & ~new_n583;
  assign new_n1768 = ~new_n583 & new_n1767;
  assign new_n1769 = ~new_n583 & ~new_n1768;
  assign new_n1770 = new_n578 & ~new_n1769;
  assign new_n1771 = new_n578 & new_n1770;
  assign new_n1772 = ~new_n1766 & ~new_n1771;
  assign new_n1773 = ~new_n662 & ~new_n1772;
  assign new_n1774 = new_n661 & new_n1773;
  assign new_n1775 = \V32(8)  & new_n662;
  assign new_n1776 = ~new_n661 & new_n1775;
  assign \V1213(8)  = new_n1774 | new_n1776;
  assign V545 = new_n538 & \V1213(8) ;
  assign new_n1779 = \V257(4)  & ~new_n534;
  assign new_n1780 = ~new_n542 & new_n1779;
  assign new_n1781 = new_n557 & new_n1780;
  assign new_n1782 = \V229(3)  & ~new_n545;
  assign new_n1783 = new_n567 & new_n1782;
  assign new_n1784 = \V189(3)  & new_n545;
  assign new_n1785 = ~new_n567 & new_n1784;
  assign new_n1786 = ~new_n1783 & ~new_n1785;
  assign new_n1787 = new_n534 & ~new_n1786;
  assign new_n1788 = ~new_n542 & new_n1787;
  assign new_n1789 = ~new_n557 & new_n1788;
  assign new_n1790 = ~new_n1781 & ~new_n1789;
  assign new_n1791 = ~new_n578 & ~new_n1790;
  assign new_n1792 = ~new_n578 & new_n1791;
  assign new_n1793 = \V32(2)  & ~new_n583;
  assign new_n1794 = ~new_n583 & new_n1793;
  assign new_n1795 = ~new_n583 & ~new_n1794;
  assign new_n1796 = new_n578 & ~new_n1795;
  assign new_n1797 = new_n578 & new_n1796;
  assign new_n1798 = ~new_n1792 & ~new_n1797;
  assign new_n1799 = ~new_n662 & ~new_n1798;
  assign new_n1800 = new_n661 & new_n1799;
  assign new_n1801 = \V32(9)  & new_n662;
  assign new_n1802 = ~new_n661 & new_n1801;
  assign \V1213(9)  = new_n1800 | new_n1802;
  assign V546 = new_n538 & \V1213(9) ;
  assign new_n1805 = \V257(5)  & ~new_n534;
  assign new_n1806 = ~new_n542 & new_n1805;
  assign new_n1807 = new_n557 & new_n1806;
  assign new_n1808 = \V229(4)  & ~new_n545;
  assign new_n1809 = new_n567 & new_n1808;
  assign new_n1810 = \V189(4)  & new_n545;
  assign new_n1811 = ~new_n567 & new_n1810;
  assign new_n1812 = ~new_n1809 & ~new_n1811;
  assign new_n1813 = new_n534 & ~new_n1812;
  assign new_n1814 = ~new_n542 & new_n1813;
  assign new_n1815 = ~new_n557 & new_n1814;
  assign new_n1816 = ~new_n1807 & ~new_n1815;
  assign new_n1817 = ~new_n578 & ~new_n1816;
  assign new_n1818 = ~new_n578 & new_n1817;
  assign new_n1819 = \V32(0)  & new_n583;
  assign new_n1820 = \V32(3)  & ~new_n583;
  assign new_n1821 = ~new_n583 & new_n1820;
  assign new_n1822 = ~new_n1819 & ~new_n1821;
  assign new_n1823 = new_n578 & ~new_n1822;
  assign new_n1824 = new_n578 & new_n1823;
  assign new_n1825 = ~new_n1818 & ~new_n1824;
  assign new_n1826 = ~new_n662 & ~new_n1825;
  assign new_n1827 = new_n661 & new_n1826;
  assign new_n1828 = \V32(10)  & new_n662;
  assign new_n1829 = ~new_n661 & new_n1828;
  assign \V1213(10)  = new_n1827 | new_n1829;
  assign V547 = new_n538 & \V1213(10) ;
  assign new_n1832 = \V229(5)  & ~new_n545;
  assign new_n1833 = new_n567 & new_n1832;
  assign new_n1834 = \V189(5)  & new_n545;
  assign new_n1835 = ~new_n567 & new_n1834;
  assign new_n1836 = ~new_n1833 & ~new_n1835;
  assign new_n1837 = new_n534 & ~new_n1836;
  assign new_n1838 = ~new_n542 & new_n1837;
  assign new_n1839 = ~new_n557 & new_n1838;
  assign new_n1840 = ~new_n1663 & ~new_n1839;
  assign new_n1841 = ~new_n578 & ~new_n1840;
  assign new_n1842 = ~new_n578 & new_n1841;
  assign new_n1843 = \V32(1)  & new_n583;
  assign new_n1844 = \V32(4)  & ~new_n583;
  assign new_n1845 = ~new_n583 & new_n1844;
  assign new_n1846 = ~new_n1843 & ~new_n1845;
  assign new_n1847 = new_n578 & ~new_n1846;
  assign new_n1848 = new_n578 & new_n1847;
  assign new_n1849 = ~new_n1842 & ~new_n1848;
  assign new_n1850 = ~new_n662 & ~new_n1849;
  assign new_n1851 = new_n661 & new_n1850;
  assign new_n1852 = \V32(11)  & new_n662;
  assign new_n1853 = ~new_n661 & new_n1852;
  assign \V1213(11)  = new_n1851 | new_n1853;
  assign V548 = new_n538 & \V1213(11) ;
  assign new_n1856 = ~\V802(0)  & ~new_n540;
  assign new_n1857 = ~new_n567 & new_n1856;
  assign new_n1858 = \V194(0)  & new_n1414;
  assign new_n1859 = \V271(0)  & ~new_n598;
  assign new_n1860 = ~\V274(0)  & new_n1859;
  assign new_n1861 = ~new_n1858 & new_n1860;
  assign new_n1862 = new_n540 & new_n1861;
  assign new_n1863 = \V134(0)  & new_n1862;
  assign new_n1864 = \V134(1)  & new_n1863;
  assign new_n1865 = ~new_n1857 & ~new_n1864;
  assign new_n1866 = \V802(0)  & new_n537;
  assign new_n1867 = \V802(0)  & \V1243(9) ;
  assign new_n1868 = new_n538 & new_n1867;
  assign new_n1869 = new_n1865 & new_n1868;
  assign new_n1870 = ~new_n1866 & new_n1869;
  assign new_n1871 = \V802(0)  & new_n538;
  assign new_n1872 = ~\V199(4)  & ~new_n1866;
  assign new_n1873 = ~new_n1865 & new_n1872;
  assign new_n1874 = ~new_n1871 & new_n1873;
  assign \V572(9)  = new_n1870 | new_n1874;
  assign new_n1876 = \V802(0)  & \V1243(8) ;
  assign new_n1877 = new_n538 & new_n1876;
  assign new_n1878 = new_n1865 & new_n1877;
  assign new_n1879 = ~new_n1866 & new_n1878;
  assign new_n1880 = ~\V199(4)  & \V199(3) ;
  assign new_n1881 = \V199(4)  & ~\V199(3) ;
  assign new_n1882 = ~new_n1880 & ~new_n1881;
  assign new_n1883 = ~new_n1866 & ~new_n1882;
  assign new_n1884 = ~new_n1865 & new_n1883;
  assign new_n1885 = ~new_n1871 & new_n1884;
  assign \V572(8)  = new_n1879 | new_n1885;
  assign new_n1887 = \V802(0)  & \V1243(7) ;
  assign new_n1888 = new_n538 & new_n1887;
  assign new_n1889 = new_n1865 & new_n1888;
  assign new_n1890 = ~new_n1866 & new_n1889;
  assign new_n1891 = \V199(4)  & \V199(3) ;
  assign new_n1892 = \V199(2)  & ~new_n1891;
  assign new_n1893 = ~\V199(2)  & new_n1891;
  assign new_n1894 = ~new_n1892 & ~new_n1893;
  assign new_n1895 = ~new_n1866 & ~new_n1894;
  assign new_n1896 = ~new_n1865 & new_n1895;
  assign new_n1897 = ~new_n1871 & new_n1896;
  assign \V572(7)  = new_n1890 | new_n1897;
  assign new_n1899 = \V239(1)  & ~new_n545;
  assign new_n1900 = new_n567 & new_n1899;
  assign new_n1901 = \V199(1)  & new_n545;
  assign new_n1902 = ~new_n567 & new_n1901;
  assign new_n1903 = ~new_n1900 & ~new_n1902;
  assign new_n1904 = ~new_n557 & ~new_n1903;
  assign new_n1905 = new_n534 & new_n1904;
  assign new_n1906 = ~new_n542 & new_n1905;
  assign new_n1907 = ~new_n578 & new_n1906;
  assign new_n1908 = ~new_n578 & new_n1907;
  assign new_n1909 = \V32(8)  & new_n583;
  assign new_n1910 = \V32(11)  & ~new_n583;
  assign new_n1911 = ~new_n583 & new_n1910;
  assign new_n1912 = ~new_n1909 & ~new_n1911;
  assign new_n1913 = new_n578 & ~new_n1912;
  assign new_n1914 = new_n578 & new_n1913;
  assign new_n1915 = ~new_n1908 & ~new_n1914;
  assign new_n1916 = ~new_n662 & ~new_n1915;
  assign new_n1917 = new_n661 & new_n1916;
  assign new_n1918 = \V84(4)  & new_n662;
  assign new_n1919 = ~new_n661 & new_n1918;
  assign \V1243(6)  = new_n1917 | new_n1919;
  assign new_n1921 = \V802(0)  & \V1243(6) ;
  assign new_n1922 = new_n538 & new_n1921;
  assign new_n1923 = new_n1865 & new_n1922;
  assign new_n1924 = ~new_n1866 & new_n1923;
  assign new_n1925 = \V199(3)  & new_n1407;
  assign new_n1926 = \V199(1)  & ~new_n1925;
  assign new_n1927 = ~\V199(1)  & new_n1925;
  assign new_n1928 = ~new_n1926 & ~new_n1927;
  assign new_n1929 = ~new_n1866 & ~new_n1928;
  assign new_n1930 = ~new_n1865 & new_n1929;
  assign new_n1931 = ~new_n1871 & new_n1930;
  assign \V572(6)  = new_n1924 | new_n1931;
  assign new_n1933 = \V239(0)  & ~new_n545;
  assign new_n1934 = new_n567 & new_n1933;
  assign new_n1935 = \V199(0)  & new_n545;
  assign new_n1936 = ~new_n567 & new_n1935;
  assign new_n1937 = ~new_n1934 & ~new_n1936;
  assign new_n1938 = ~new_n557 & ~new_n1937;
  assign new_n1939 = new_n534 & new_n1938;
  assign new_n1940 = ~new_n542 & new_n1939;
  assign new_n1941 = ~new_n578 & new_n1940;
  assign new_n1942 = ~new_n578 & new_n1941;
  assign new_n1943 = \V32(7)  & new_n583;
  assign new_n1944 = \V32(10)  & ~new_n583;
  assign new_n1945 = ~new_n583 & new_n1944;
  assign new_n1946 = ~new_n1943 & ~new_n1945;
  assign new_n1947 = new_n578 & ~new_n1946;
  assign new_n1948 = new_n578 & new_n1947;
  assign new_n1949 = ~new_n1942 & ~new_n1948;
  assign new_n1950 = ~new_n662 & ~new_n1949;
  assign new_n1951 = new_n661 & new_n1950;
  assign new_n1952 = \V84(3)  & new_n662;
  assign new_n1953 = ~new_n661 & new_n1952;
  assign \V1243(5)  = new_n1951 | new_n1953;
  assign new_n1955 = \V802(0)  & \V1243(5) ;
  assign new_n1956 = new_n538 & new_n1955;
  assign new_n1957 = new_n1865 & new_n1956;
  assign new_n1958 = ~new_n1866 & new_n1957;
  assign new_n1959 = \V199(1)  & new_n1407;
  assign new_n1960 = \V199(3)  & new_n1959;
  assign new_n1961 = \V199(0)  & ~new_n1960;
  assign new_n1962 = ~\V199(0)  & new_n1960;
  assign new_n1963 = ~new_n1961 & ~new_n1962;
  assign new_n1964 = ~new_n1866 & ~new_n1963;
  assign new_n1965 = ~new_n1865 & new_n1964;
  assign new_n1966 = ~new_n1871 & new_n1965;
  assign \V572(5)  = new_n1958 | new_n1966;
  assign new_n1968 = \V234(4)  & ~new_n545;
  assign new_n1969 = new_n567 & new_n1968;
  assign new_n1970 = \V194(4)  & new_n545;
  assign new_n1971 = ~new_n567 & new_n1970;
  assign new_n1972 = ~new_n1969 & ~new_n1971;
  assign new_n1973 = ~new_n557 & ~new_n1972;
  assign new_n1974 = new_n534 & new_n1973;
  assign new_n1975 = ~new_n542 & new_n1974;
  assign new_n1976 = ~new_n578 & new_n1975;
  assign new_n1977 = ~new_n578 & new_n1976;
  assign new_n1978 = \V32(6)  & new_n583;
  assign new_n1979 = \V32(9)  & ~new_n583;
  assign new_n1980 = ~new_n583 & new_n1979;
  assign new_n1981 = ~new_n1978 & ~new_n1980;
  assign new_n1982 = new_n578 & ~new_n1981;
  assign new_n1983 = new_n578 & new_n1982;
  assign new_n1984 = ~new_n1977 & ~new_n1983;
  assign new_n1985 = ~new_n662 & ~new_n1984;
  assign new_n1986 = new_n661 & new_n1985;
  assign new_n1987 = \V84(2)  & new_n662;
  assign new_n1988 = ~new_n661 & new_n1987;
  assign \V1243(4)  = new_n1986 | new_n1988;
  assign new_n1990 = \V802(0)  & \V1243(4) ;
  assign new_n1991 = new_n538 & new_n1990;
  assign new_n1992 = new_n1865 & new_n1991;
  assign new_n1993 = ~new_n1866 & new_n1992;
  assign new_n1994 = \V199(1)  & new_n1408;
  assign new_n1995 = \V199(3)  & new_n1994;
  assign new_n1996 = \V194(4)  & ~new_n1995;
  assign new_n1997 = ~\V194(4)  & new_n1995;
  assign new_n1998 = ~new_n1996 & ~new_n1997;
  assign new_n1999 = ~new_n1866 & ~new_n1998;
  assign new_n2000 = ~new_n1865 & new_n1999;
  assign new_n2001 = ~new_n1871 & new_n2000;
  assign \V572(4)  = new_n1993 | new_n2001;
  assign new_n2003 = \V149(7)  & \V802(0) ;
  assign new_n2004 = new_n537 & new_n2003;
  assign new_n2005 = new_n1865 & new_n2004;
  assign new_n2006 = ~new_n1871 & new_n2005;
  assign new_n2007 = \V194(4)  & new_n1408;
  assign new_n2008 = \V199(1)  & new_n2007;
  assign new_n2009 = \V199(3)  & new_n2008;
  assign new_n2010 = \V194(3)  & ~new_n2009;
  assign new_n2011 = ~\V194(3)  & new_n2009;
  assign new_n2012 = ~new_n2010 & ~new_n2011;
  assign new_n2013 = ~new_n1866 & ~new_n2012;
  assign new_n2014 = ~new_n1865 & new_n2013;
  assign new_n2015 = ~new_n1871 & new_n2014;
  assign new_n2016 = \V234(3)  & ~new_n545;
  assign new_n2017 = new_n567 & new_n2016;
  assign new_n2018 = \V194(3)  & new_n545;
  assign new_n2019 = ~new_n567 & new_n2018;
  assign new_n2020 = ~new_n2017 & ~new_n2019;
  assign new_n2021 = new_n534 & ~new_n2020;
  assign new_n2022 = ~new_n542 & new_n2021;
  assign new_n2023 = ~new_n557 & new_n2022;
  assign new_n2024 = ~\V59(0)  & \V149(7) ;
  assign new_n2025 = ~new_n540 & new_n2024;
  assign new_n2026 = new_n537 & new_n2025;
  assign new_n2027 = new_n534 & new_n2026;
  assign new_n2028 = new_n557 & new_n2027;
  assign new_n2029 = ~new_n2023 & ~new_n2028;
  assign new_n2030 = ~new_n578 & ~new_n2029;
  assign new_n2031 = ~new_n578 & new_n2030;
  assign new_n2032 = \V32(5)  & new_n583;
  assign new_n2033 = \V32(8)  & ~new_n583;
  assign new_n2034 = ~new_n583 & new_n2033;
  assign new_n2035 = ~new_n2032 & ~new_n2034;
  assign new_n2036 = new_n578 & ~new_n2035;
  assign new_n2037 = new_n578 & new_n2036;
  assign new_n2038 = ~new_n2031 & ~new_n2037;
  assign new_n2039 = ~new_n662 & ~new_n2038;
  assign new_n2040 = new_n661 & new_n2039;
  assign new_n2041 = \V84(1)  & new_n662;
  assign new_n2042 = ~new_n661 & new_n2041;
  assign \V1243(3)  = new_n2040 | new_n2042;
  assign new_n2044 = \V802(0)  & \V1243(3) ;
  assign new_n2045 = new_n538 & new_n2044;
  assign new_n2046 = new_n1865 & new_n2045;
  assign new_n2047 = ~new_n1866 & new_n2046;
  assign new_n2048 = ~new_n2006 & ~new_n2015;
  assign \V572(3)  = new_n2047 | ~new_n2048;
  assign new_n2050 = \V149(6)  & \V802(0) ;
  assign new_n2051 = new_n537 & new_n2050;
  assign new_n2052 = new_n1865 & new_n2051;
  assign new_n2053 = ~new_n1871 & new_n2052;
  assign new_n2054 = \V194(4)  & new_n1409;
  assign new_n2055 = \V199(1)  & new_n2054;
  assign new_n2056 = \V199(3)  & new_n2055;
  assign new_n2057 = \V194(2)  & ~new_n2056;
  assign new_n2058 = ~\V194(2)  & new_n2056;
  assign new_n2059 = ~new_n2057 & ~new_n2058;
  assign new_n2060 = ~new_n1866 & ~new_n2059;
  assign new_n2061 = ~new_n1865 & new_n2060;
  assign new_n2062 = ~new_n1871 & new_n2061;
  assign new_n2063 = \V234(2)  & ~new_n545;
  assign new_n2064 = new_n567 & new_n2063;
  assign new_n2065 = \V194(2)  & new_n545;
  assign new_n2066 = ~new_n567 & new_n2065;
  assign new_n2067 = ~new_n2064 & ~new_n2066;
  assign new_n2068 = new_n534 & ~new_n2067;
  assign new_n2069 = ~new_n542 & new_n2068;
  assign new_n2070 = ~new_n557 & new_n2069;
  assign new_n2071 = ~\V59(0)  & \V149(6) ;
  assign new_n2072 = ~new_n540 & new_n2071;
  assign new_n2073 = new_n537 & new_n2072;
  assign new_n2074 = new_n534 & new_n2073;
  assign new_n2075 = new_n557 & new_n2074;
  assign new_n2076 = ~new_n2070 & ~new_n2075;
  assign new_n2077 = ~new_n578 & ~new_n2076;
  assign new_n2078 = ~new_n578 & new_n2077;
  assign new_n2079 = \V32(4)  & new_n583;
  assign new_n2080 = \V32(7)  & ~new_n583;
  assign new_n2081 = ~new_n583 & new_n2080;
  assign new_n2082 = ~new_n2079 & ~new_n2081;
  assign new_n2083 = new_n578 & ~new_n2082;
  assign new_n2084 = new_n578 & new_n2083;
  assign new_n2085 = ~new_n2078 & ~new_n2084;
  assign new_n2086 = ~new_n662 & ~new_n2085;
  assign new_n2087 = new_n661 & new_n2086;
  assign new_n2088 = \V84(0)  & new_n662;
  assign new_n2089 = ~new_n661 & new_n2088;
  assign \V1243(2)  = new_n2087 | new_n2089;
  assign new_n2091 = \V802(0)  & \V1243(2) ;
  assign new_n2092 = new_n538 & new_n2091;
  assign new_n2093 = new_n1865 & new_n2092;
  assign new_n2094 = ~new_n1866 & new_n2093;
  assign new_n2095 = ~new_n2053 & ~new_n2062;
  assign \V572(2)  = new_n2094 | ~new_n2095;
  assign new_n2097 = \V149(5)  & \V802(0) ;
  assign new_n2098 = new_n537 & new_n2097;
  assign new_n2099 = new_n1865 & new_n2098;
  assign new_n2100 = ~new_n1871 & new_n2099;
  assign new_n2101 = \V194(2)  & new_n1409;
  assign new_n2102 = \V194(4)  & new_n2101;
  assign new_n2103 = \V199(1)  & new_n2102;
  assign new_n2104 = \V199(3)  & new_n2103;
  assign new_n2105 = \V194(1)  & ~new_n2104;
  assign new_n2106 = ~\V194(1)  & new_n2104;
  assign new_n2107 = ~new_n2105 & ~new_n2106;
  assign new_n2108 = ~new_n1866 & ~new_n2107;
  assign new_n2109 = ~new_n1865 & new_n2108;
  assign new_n2110 = ~new_n1871 & new_n2109;
  assign new_n2111 = \V234(1)  & ~new_n545;
  assign new_n2112 = new_n567 & new_n2111;
  assign new_n2113 = \V194(1)  & new_n545;
  assign new_n2114 = ~new_n567 & new_n2113;
  assign new_n2115 = ~new_n2112 & ~new_n2114;
  assign new_n2116 = new_n534 & ~new_n2115;
  assign new_n2117 = ~new_n542 & new_n2116;
  assign new_n2118 = ~new_n557 & new_n2117;
  assign new_n2119 = ~\V59(0)  & \V149(5) ;
  assign new_n2120 = ~new_n540 & new_n2119;
  assign new_n2121 = new_n537 & new_n2120;
  assign new_n2122 = new_n534 & new_n2121;
  assign new_n2123 = new_n557 & new_n2122;
  assign new_n2124 = ~new_n2118 & ~new_n2123;
  assign new_n2125 = ~new_n578 & ~new_n2124;
  assign new_n2126 = ~new_n578 & new_n2125;
  assign new_n2127 = \V32(3)  & new_n583;
  assign new_n2128 = \V32(6)  & ~new_n583;
  assign new_n2129 = ~new_n583 & new_n2128;
  assign new_n2130 = ~new_n2127 & ~new_n2129;
  assign new_n2131 = new_n578 & ~new_n2130;
  assign new_n2132 = new_n578 & new_n2131;
  assign new_n2133 = ~new_n2126 & ~new_n2132;
  assign new_n2134 = ~new_n662 & ~new_n2133;
  assign new_n2135 = new_n661 & new_n2134;
  assign new_n2136 = \V78(5)  & new_n662;
  assign new_n2137 = ~new_n661 & new_n2136;
  assign \V1243(1)  = new_n2135 | new_n2137;
  assign new_n2139 = \V802(0)  & \V1243(1) ;
  assign new_n2140 = new_n538 & new_n2139;
  assign new_n2141 = new_n1865 & new_n2140;
  assign new_n2142 = ~new_n1866 & new_n2141;
  assign new_n2143 = ~new_n2100 & ~new_n2110;
  assign \V572(1)  = new_n2142 | ~new_n2143;
  assign new_n2145 = \V149(4)  & \V802(0) ;
  assign new_n2146 = new_n537 & new_n2145;
  assign new_n2147 = new_n1865 & new_n2146;
  assign new_n2148 = ~new_n1871 & new_n2147;
  assign new_n2149 = \V194(0)  & ~new_n1414;
  assign new_n2150 = ~\V194(0)  & new_n1414;
  assign new_n2151 = ~new_n2149 & ~new_n2150;
  assign new_n2152 = ~new_n1866 & ~new_n2151;
  assign new_n2153 = ~new_n1865 & new_n2152;
  assign new_n2154 = ~new_n1871 & new_n2153;
  assign new_n2155 = \V802(0)  & ~\V321(2) ;
  assign new_n2156 = new_n538 & new_n2155;
  assign new_n2157 = new_n1865 & new_n2156;
  assign new_n2158 = ~new_n1866 & new_n2157;
  assign new_n2159 = ~new_n2148 & ~new_n2154;
  assign \V572(0)  = new_n2158 | ~new_n2159;
  assign new_n2161 = \V802(0)  & ~new_n567;
  assign V587 = ~\V243(0)  & ~new_n2161;
  assign new_n2163 = ~\V243(0)  & \V244(0) ;
  assign new_n2164 = ~new_n2161 & new_n2163;
  assign new_n2165 = \V243(0)  & ~\V244(0) ;
  assign new_n2166 = ~new_n2161 & new_n2165;
  assign \V591(0)  = new_n2164 | new_n2166;
  assign new_n2168 = \V245(0)  & ~new_n1307;
  assign new_n2169 = ~new_n2161 & new_n2168;
  assign new_n2170 = ~\V245(0)  & new_n1307;
  assign new_n2171 = ~new_n2161 & new_n2170;
  assign \V597(0)  = new_n2169 | new_n2171;
  assign new_n2173 = \V246(0)  & ~new_n1308;
  assign new_n2174 = ~new_n2161 & new_n2173;
  assign new_n2175 = ~\V246(0)  & new_n1308;
  assign new_n2176 = ~new_n2161 & new_n2175;
  assign \V603(0)  = new_n2174 | new_n2176;
  assign new_n2178 = \V247(0)  & ~new_n1309;
  assign new_n2179 = ~new_n2161 & new_n2178;
  assign new_n2180 = ~\V247(0)  & new_n1309;
  assign new_n2181 = ~new_n2161 & new_n2180;
  assign \V609(0)  = new_n2179 | new_n2181;
  assign new_n2183 = \V62(0)  & ~\V214(0) ;
  assign new_n2184 = new_n1513 & new_n2183;
  assign new_n2185 = ~new_n1311 & new_n2184;
  assign new_n2186 = ~new_n1311 & ~new_n1586;
  assign new_n2187 = new_n1626 & new_n2186;
  assign new_n2188 = ~\V214(0)  & new_n2187;
  assign new_n2189 = ~new_n631 & ~new_n1620;
  assign new_n2190 = \V59(0)  & ~\V214(0) ;
  assign new_n2191 = ~new_n2189 & new_n2190;
  assign new_n2192 = ~new_n1311 & new_n2191;
  assign new_n2193 = ~new_n2185 & ~new_n2188;
  assign V620 = ~new_n2192 & new_n2193;
  assign new_n2195 = ~\V45(0)  & \V41(0) ;
  assign new_n2196 = \V45(0)  & ~\V41(0) ;
  assign new_n2197 = ~new_n2195 & ~new_n2196;
  assign V621 = \V293(0)  & new_n2197;
  assign new_n2199 = \V274(0)  & ~\V202(0) ;
  assign new_n2200 = ~\V271(0)  & new_n2199;
  assign \V640(0)  = \V271(0)  | new_n2200;
  assign new_n2202 = \V274(0)  & ~\V640(0) ;
  assign new_n2203 = \V271(0)  & ~new_n2200;
  assign new_n2204 = \V269(0)  & new_n2203;
  assign \V634(0)  = ~new_n2202 & ~new_n2204;
  assign new_n2206 = ~\V290(0)  & new_n1311;
  assign new_n2207 = \V165(7)  & new_n2206;
  assign new_n2208 = \V261(0)  & ~new_n1604;
  assign new_n2209 = ~\V802(0)  & new_n2208;
  assign new_n2210 = \V272(0)  & new_n2209;
  assign new_n2211 = ~\V275(0)  & new_n2210;
  assign new_n2212 = new_n540 & new_n2211;
  assign new_n2213 = ~\V149(6)  & new_n1510;
  assign new_n2214 = ~new_n544 & new_n2213;
  assign new_n2215 = new_n1586 & new_n2214;
  assign new_n2216 = \V62(0)  & new_n2215;
  assign new_n2217 = ~new_n544 & new_n627;
  assign new_n2218 = new_n1586 & new_n2217;
  assign new_n2219 = \V59(0)  & new_n2218;
  assign new_n2220 = \V67(0)  & \V172(0) ;
  assign new_n2221 = \V215(0)  & new_n2220;
  assign new_n2222 = ~new_n544 & new_n1586;
  assign new_n2223 = ~new_n1509 & new_n2222;
  assign new_n2224 = ~new_n2213 & new_n2223;
  assign new_n2225 = ~new_n627 & new_n2224;
  assign new_n2226 = \V59(0)  & ~new_n544;
  assign new_n2227 = new_n1586 & new_n2226;
  assign new_n2228 = new_n1509 & new_n2227;
  assign new_n2229 = ~new_n2221 & ~new_n2225;
  assign new_n2230 = ~new_n2228 & new_n2229;
  assign new_n2231 = ~new_n2216 & ~new_n2219;
  assign new_n2232 = ~\V214(0)  & new_n2231;
  assign new_n2233 = new_n2230 & new_n2232;
  assign new_n2234 = \V56(0)  & ~new_n566;
  assign new_n2235 = ~new_n540 & ~new_n2234;
  assign new_n2236 = \V242(0)  & new_n2235;
  assign new_n2237 = ~\V802(0)  & new_n2236;
  assign new_n2238 = ~new_n567 & new_n2237;
  assign new_n2239 = \V261(0)  & ~new_n540;
  assign new_n2240 = ~new_n1604 & new_n2239;
  assign new_n2241 = ~\V802(0)  & new_n2240;
  assign new_n2242 = \V134(1)  & \V134(0) ;
  assign new_n2243 = \V242(0)  & new_n2242;
  assign new_n2244 = ~\V802(0)  & new_n2243;
  assign new_n2245 = \V272(0)  & new_n2244;
  assign new_n2246 = ~\V275(0)  & new_n2245;
  assign new_n2247 = new_n540 & new_n2246;
  assign new_n2248 = ~new_n2241 & ~new_n2247;
  assign new_n2249 = ~new_n2212 & new_n2233;
  assign new_n2250 = ~new_n2238 & new_n2249;
  assign new_n2251 = new_n2248 & new_n2250;
  assign new_n2252 = ~new_n1457 & new_n2251;
  assign new_n2253 = ~\V302(0)  & ~new_n2207;
  assign new_n2254 = new_n2252 & new_n2253;
  assign new_n2255 = \V70(0)  & ~new_n533;
  assign new_n2256 = V763 & new_n2255;
  assign new_n2257 = new_n2254 & new_n2256;
  assign V775 = \V14(0)  & new_n2257;
  assign new_n2259 = \V10(0)  & ~\V13(0) ;
  assign V779 = \V6(0)  & new_n2259;
  assign new_n2261 = \V56(0)  & ~new_n500;
  assign new_n2262 = ~\V174(0)  & new_n2261;
  assign new_n2263 = ~\V52(0)  & ~new_n2262;
  assign new_n2264 = \V12(0)  & ~new_n2263;
  assign V781 = \V6(0)  & new_n2264;
  assign V782 = \V7(0)  & new_n2259;
  assign V783 = \V5(0)  & \V11(0) ;
  assign V784 = \V7(0)  & \V11(0) ;
  assign new_n2269 = ~\V149(7)  & ~\V149(3) ;
  assign new_n2270 = \V149(4)  & new_n2269;
  assign new_n2271 = new_n489 & new_n2270;
  assign new_n2272 = \V149(5)  & new_n2271;
  assign new_n2273 = ~\V149(6)  & new_n2272;
  assign new_n2274 = \V149(3)  & new_n594;
  assign new_n2275 = new_n489 & new_n2274;
  assign new_n2276 = ~\V149(4)  & new_n2275;
  assign new_n2277 = ~\V149(6)  & new_n2276;
  assign new_n2278 = \V149(6)  & new_n671;
  assign new_n2279 = ~new_n672 & ~new_n2277;
  assign new_n2280 = new_n489 & new_n2279;
  assign new_n2281 = \V149(3)  & new_n2280;
  assign new_n2282 = ~new_n2278 & new_n2281;
  assign new_n2283 = ~\V149(4)  & new_n1574;
  assign new_n2284 = ~\V149(6)  & new_n2283;
  assign new_n2285 = ~new_n2273 & ~new_n2282;
  assign new_n2286 = ~new_n2284 & new_n2285;
  assign new_n2287 = ~\V302(0)  & ~new_n2286;
  assign new_n2288 = \V149(0)  & \V149(2) ;
  assign new_n2289 = \V149(1)  & new_n2288;
  assign new_n2290 = \V149(0)  & ~\V149(1) ;
  assign new_n2291 = \V149(2)  & new_n2290;
  assign new_n2292 = \V149(0)  & ~\V149(2) ;
  assign new_n2293 = \V149(1)  & new_n2292;
  assign new_n2294 = ~new_n2289 & ~new_n2291;
  assign new_n2295 = new_n2286 & new_n2294;
  assign new_n2296 = ~new_n2293 & new_n2295;
  assign new_n2297 = new_n534 & ~new_n2287;
  assign new_n2298 = ~new_n2296 & new_n2297;
  assign new_n2299 = \V290(0)  & ~new_n1311;
  assign new_n2300 = ~\V149(6)  & new_n493;
  assign new_n2301 = ~\V149(6)  & new_n1575;
  assign new_n2302 = ~\V59(0)  & ~new_n534;
  assign new_n2303 = ~\V259(0)  & new_n2302;
  assign new_n2304 = ~\V260(0)  & new_n2303;
  assign new_n2305 = \V258(0)  & new_n2304;
  assign new_n2306 = \V149(6)  & new_n2283;
  assign new_n2307 = ~\V149(6)  & new_n597;
  assign new_n2308 = ~\V149(6)  & new_n1502;
  assign new_n2309 = ~new_n1576 & ~new_n2300;
  assign new_n2310 = ~new_n2301 & new_n2309;
  assign new_n2311 = ~new_n2305 & new_n2310;
  assign new_n2312 = ~new_n2306 & new_n2311;
  assign new_n2313 = ~new_n2307 & new_n2312;
  assign new_n2314 = ~new_n2308 & new_n2313;
  assign new_n2315 = \V56(0)  & ~new_n2314;
  assign new_n2316 = \V65(0)  & new_n1513;
  assign new_n2317 = ~new_n1511 & ~new_n1514;
  assign new_n2318 = \V62(0)  & ~new_n2317;
  assign new_n2319 = ~new_n2315 & ~new_n2316;
  assign new_n2320 = ~new_n2318 & new_n2319;
  assign new_n2321 = ~new_n1311 & new_n2219;
  assign new_n2322 = \V290(0)  & new_n1311;
  assign new_n2323 = ~new_n1311 & new_n2225;
  assign new_n2324 = ~new_n1311 & new_n2228;
  assign new_n2325 = ~new_n2323 & ~new_n2324;
  assign new_n2326 = ~new_n2216 & ~new_n2321;
  assign new_n2327 = ~new_n2322 & new_n2326;
  assign \V1741(0)  = ~new_n2325 | ~new_n2327;
  assign new_n2329 = ~new_n1457 & ~new_n2320;
  assign new_n2330 = ~\V1741(0)  & new_n2329;
  assign new_n2331 = ~new_n1304 & new_n2254;
  assign new_n2332 = ~new_n1604 & ~new_n2331;
  assign new_n2333 = ~\V289(0)  & ~new_n2330;
  assign new_n2334 = ~\V302(0)  & ~new_n2299;
  assign new_n2335 = new_n2333 & new_n2334;
  assign new_n2336 = ~\V214(0)  & ~new_n2332;
  assign new_n2337 = ~new_n2207 & new_n2336;
  assign new_n2338 = new_n2335 & new_n2337;
  assign new_n2339 = \V14(0)  & ~new_n2298;
  assign \V798(0)  = ~new_n2338 | ~new_n2339;
  assign V801 = new_n500 & new_n509;
  assign new_n2342 = \V802(0)  & new_n591;
  assign new_n2343 = ~\V279(0)  & ~new_n2342;
  assign new_n2344 = \V149(5)  & new_n2342;
  assign \V821(0)  = new_n2343 | new_n2344;
  assign new_n2346 = \V280(0)  & ~new_n2342;
  assign new_n2347 = \V279(0)  & new_n2346;
  assign new_n2348 = \V149(4)  & new_n2342;
  assign new_n2349 = ~\V280(0)  & new_n2343;
  assign new_n2350 = ~new_n2347 & ~new_n2348;
  assign \V826(0)  = new_n2349 | ~new_n2350;
  assign new_n2352 = ~new_n500 & new_n509;
  assign new_n2353 = \V56(0)  & V763;
  assign new_n2354 = ~new_n500 & new_n2353;
  assign new_n2355 = ~new_n2263 & new_n2354;
  assign new_n2356 = \V802(0)  & ~new_n2298;
  assign new_n2357 = \V56(0)  & ~new_n2286;
  assign new_n2358 = ~new_n2356 & ~new_n2357;
  assign new_n2359 = ~new_n2352 & ~new_n2355;
  assign new_n2360 = new_n2358 & new_n2359;
  assign new_n2361 = new_n2254 & ~new_n2360;
  assign V966 = \V14(0)  & new_n2361;
  assign new_n2363 = \V62(0)  & ~new_n534;
  assign new_n2364 = \V56(0)  & new_n2286;
  assign new_n2365 = new_n2314 & new_n2364;
  assign new_n2366 = ~new_n2355 & new_n2365;
  assign new_n2367 = new_n567 & ~new_n591;
  assign new_n2368 = ~new_n1621 & new_n2367;
  assign new_n2369 = \V59(0)  & ~new_n2368;
  assign new_n2370 = ~new_n2363 & ~new_n2366;
  assign new_n2371 = ~new_n2369 & new_n2370;
  assign new_n2372 = new_n2254 & ~new_n2371;
  assign V986 = \V14(0)  & new_n2372;
  assign V1256 = \V2(0)  & new_n2259;
  assign new_n2375 = ~\V57(0)  & new_n1514;
  assign new_n2376 = ~new_n630 & new_n647;
  assign new_n2377 = ~new_n538 & new_n2376;
  assign new_n2378 = ~new_n591 & new_n1429;
  assign new_n2379 = new_n626 & new_n2378;
  assign new_n2380 = new_n2377 & new_n2379;
  assign new_n2381 = \V57(0)  & ~new_n2380;
  assign new_n2382 = ~\V60(0)  & ~\V63(0) ;
  assign new_n2383 = new_n598 & ~new_n2382;
  assign new_n2384 = \V12(0)  & \V2(0) ;
  assign new_n2385 = ~\V174(0)  & new_n2384;
  assign new_n2386 = ~new_n2375 & new_n2385;
  assign new_n2387 = ~new_n2381 & new_n2386;
  assign new_n2388 = ~new_n2383 & new_n2387;
  assign V1257 = ~\V35(0)  & new_n2388;
  assign V1260 = \V11(0)  & \V3(0) ;
  assign V1261 = ~\V62(0)  & V1260;
  assign V1262 = \V4(0)  & new_n2259;
  assign V1264 = \V12(0)  & \V4(0) ;
  assign V1265 = \V52(0)  & V1264;
  assign V1266 = \V11(0)  & \V4(0) ;
  assign V1267 = \V11(0)  & \V2(0) ;
  assign new_n2397 = \V14(0)  & new_n2254;
  assign new_n2398 = new_n631 & new_n2397;
  assign new_n2399 = \V62(0)  & new_n2398;
  assign new_n2400 = ~new_n538 & ~new_n1621;
  assign new_n2401 = ~new_n537 & ~new_n1426;
  assign new_n2402 = new_n2400 & new_n2401;
  assign new_n2403 = ~new_n549 & ~new_n1430;
  assign new_n2404 = ~new_n591 & new_n2403;
  assign new_n2405 = new_n2402 & new_n2404;
  assign new_n2406 = ~\V174(0)  & new_n499;
  assign new_n2407 = \V59(0)  & ~V1719;
  assign new_n2408 = ~new_n1509 & new_n2407;
  assign new_n2409 = new_n2405 & new_n2408;
  assign new_n2410 = ~new_n2406 & new_n2409;
  assign new_n2411 = ~new_n672 & new_n2410;
  assign new_n2412 = new_n2254 & new_n2411;
  assign new_n2413 = \V14(0)  & new_n2412;
  assign \V1274(0)  = new_n2399 | new_n2413;
  assign new_n2415 = \V56(0)  & new_n2308;
  assign new_n2416 = ~\V302(0)  & new_n544;
  assign new_n2417 = new_n599 & new_n627;
  assign new_n2418 = ~new_n2213 & ~new_n2417;
  assign new_n2419 = ~new_n1509 & ~new_n2416;
  assign new_n2420 = new_n2418 & new_n2419;
  assign new_n2421 = ~\V289(0)  & \V14(0) ;
  assign new_n2422 = ~new_n2420 & new_n2421;
  assign new_n2423 = new_n1586 & new_n2422;
  assign new_n2424 = ~new_n1311 & new_n2423;
  assign new_n2425 = new_n485 & ~new_n1311;
  assign new_n2426 = new_n1586 & new_n2425;
  assign new_n2427 = ~new_n2424 & new_n2426;
  assign new_n2428 = ~new_n499 & new_n2427;
  assign new_n2429 = new_n485 & new_n2322;
  assign new_n2430 = ~new_n2428 & ~new_n2429;
  assign new_n2431 = \V14(0)  & ~new_n2415;
  assign new_n2432 = \V213(0)  & new_n2431;
  assign new_n2433 = new_n2430 & new_n2432;
  assign new_n2434 = new_n2430 & new_n2433;
  assign new_n2435 = ~\V165(5)  & ~\V165(7) ;
  assign new_n2436 = ~\V165(3)  & new_n2435;
  assign new_n2437 = ~\V165(4)  & new_n2436;
  assign new_n2438 = ~\V165(6)  & new_n2437;
  assign new_n2439 = ~new_n1586 & ~new_n2438;
  assign new_n2440 = ~new_n2430 & ~new_n2439;
  assign new_n2441 = ~new_n2430 & new_n2440;
  assign \V1281(0)  = new_n2434 | new_n2441;
  assign new_n2443 = \V213(5)  & new_n2431;
  assign new_n2444 = ~new_n2429 & new_n2443;
  assign new_n2445 = ~new_n2429 & new_n2444;
  assign new_n2446 = \V165(7)  & new_n2429;
  assign new_n2447 = new_n2429 & new_n2446;
  assign \V1297(4)  = new_n2445 | new_n2447;
  assign new_n2449 = \V213(4)  & new_n2431;
  assign new_n2450 = ~new_n2429 & new_n2449;
  assign new_n2451 = ~new_n2429 & new_n2450;
  assign new_n2452 = \V165(6)  & new_n2429;
  assign new_n2453 = new_n2429 & new_n2452;
  assign \V1297(3)  = new_n2451 | new_n2453;
  assign new_n2455 = \V213(3)  & new_n2431;
  assign new_n2456 = ~new_n2429 & new_n2455;
  assign new_n2457 = ~new_n2429 & new_n2456;
  assign new_n2458 = \V165(5)  & new_n2429;
  assign new_n2459 = new_n2429 & new_n2458;
  assign \V1297(2)  = new_n2457 | new_n2459;
  assign new_n2461 = \V213(2)  & new_n2431;
  assign new_n2462 = ~new_n2429 & new_n2461;
  assign new_n2463 = ~new_n2429 & new_n2462;
  assign new_n2464 = \V165(4)  & new_n2429;
  assign new_n2465 = new_n2429 & new_n2464;
  assign \V1297(1)  = new_n2463 | new_n2465;
  assign new_n2467 = \V213(1)  & new_n2431;
  assign new_n2468 = ~new_n2429 & new_n2467;
  assign new_n2469 = ~new_n2429 & new_n2468;
  assign new_n2470 = \V165(3)  & new_n2429;
  assign new_n2471 = new_n2429 & new_n2470;
  assign \V1297(0)  = new_n2469 | new_n2471;
  assign new_n2473 = ~new_n1514 & new_n2397;
  assign new_n2474 = ~new_n2213 & new_n2473;
  assign new_n2475 = ~new_n1440 & new_n2474;
  assign new_n2476 = new_n534 & new_n2475;
  assign new_n2477 = ~new_n1441 & new_n2476;
  assign new_n2478 = new_n647 & new_n2477;
  assign new_n2479 = ~new_n1511 & new_n2478;
  assign V1365 = \V62(0)  & new_n2479;
  assign new_n2481 = \V802(0)  & ~new_n566;
  assign V1378 = V782 & new_n2481;
  assign new_n2483 = ~\V802(0)  & new_n1858;
  assign new_n2484 = ~\V802(0)  & new_n540;
  assign new_n2485 = \V248(0)  & ~\V802(0) ;
  assign new_n2486 = ~new_n2241 & ~new_n2483;
  assign new_n2487 = ~new_n566 & new_n2486;
  assign new_n2488 = ~new_n2484 & new_n2487;
  assign new_n2489 = ~new_n2485 & new_n2488;
  assign new_n2490 = ~new_n2241 & ~new_n2485;
  assign new_n2491 = ~new_n540 & new_n2490;
  assign new_n2492 = ~\V802(0)  & new_n2491;
  assign new_n2493 = new_n549 & new_n2492;
  assign new_n2494 = ~new_n1858 & new_n2493;
  assign new_n2495 = ~new_n1864 & ~new_n2489;
  assign new_n2496 = ~new_n2494 & new_n2495;
  assign V1380 = V782 & ~new_n2496;
  assign new_n2498 = \V802(0)  & ~new_n1580;
  assign new_n2499 = ~new_n591 & ~new_n2498;
  assign new_n2500 = \V7(0)  & ~new_n2499;
  assign V1382 = new_n2259 & new_n2500;
  assign new_n2502 = \V56(0)  & ~new_n1311;
  assign new_n2503 = new_n1576 & new_n2502;
  assign new_n2504 = ~new_n1584 & new_n2503;
  assign new_n2505 = \V7(0)  & new_n2504;
  assign V1384 = new_n2259 & new_n2505;
  assign new_n2507 = ~\V56(0)  & ~\V50(0) ;
  assign new_n2508 = ~\V62(0)  & new_n2507;
  assign new_n2509 = ~new_n534 & ~new_n2508;
  assign new_n2510 = \V7(0)  & new_n2509;
  assign V1386 = new_n2259 & new_n2510;
  assign new_n2512 = V763 & new_n2397;
  assign new_n2513 = ~\V165(5)  & new_n2512;
  assign new_n2514 = \V165(3)  & new_n2513;
  assign new_n2515 = ~\V165(4)  & new_n2514;
  assign new_n2516 = \V165(6)  & new_n2515;
  assign new_n2517 = \V70(0)  & new_n2516;
  assign new_n2518 = ~new_n1513 & new_n2397;
  assign new_n2519 = \V65(0)  & new_n2518;
  assign new_n2520 = ~new_n628 & new_n2519;
  assign \V1392(0)  = new_n2517 | new_n2520;
  assign V1426 = \V1(0)  & new_n2259;
  assign V1428 = \V1(0)  & \V11(0) ;
  assign V1429 = \V1(0)  & \V12(0) ;
  assign new_n2525 = \V66(0)  & new_n2254;
  assign V1432 = \V14(0)  & new_n2525;
  assign new_n2527 = \V277(0)  & ~new_n538;
  assign new_n2528 = \V14(0)  & new_n2527;
  assign \V1439(0)  = new_n2300 | new_n2528;
  assign \V1440(0)  = ~\V14(0)  | new_n540;
  assign new_n2531 = \V268(5)  & \V268(3) ;
  assign new_n2532 = \V268(1)  & new_n2531;
  assign new_n2533 = \V268(2)  & new_n2532;
  assign new_n2534 = \V268(4)  & new_n2533;
  assign new_n2535 = \V268(0)  & new_n2534;
  assign new_n2536 = ~new_n2509 & ~new_n2535;
  assign new_n2537 = \V14(0)  & new_n2536;
  assign new_n2538 = \V258(0)  & new_n2537;
  assign new_n2539 = \V14(0)  & ~new_n2536;
  assign new_n2540 = ~\V258(0)  & new_n2539;
  assign \V1451(0)  = new_n2538 | new_n2540;
  assign new_n2542 = ~\V258(0)  & new_n2509;
  assign new_n2543 = \V258(0)  & new_n2535;
  assign new_n2544 = ~new_n2542 & ~new_n2543;
  assign new_n2545 = \V259(0)  & new_n2544;
  assign new_n2546 = \V14(0)  & new_n2545;
  assign new_n2547 = ~\V259(0)  & ~new_n2544;
  assign new_n2548 = \V14(0)  & new_n2547;
  assign \V1459(0)  = new_n2546 | new_n2548;
  assign new_n2550 = ~\V259(0)  & new_n2542;
  assign new_n2551 = \V259(0)  & new_n2543;
  assign new_n2552 = ~new_n2550 & ~new_n2551;
  assign new_n2553 = \V260(0)  & new_n2552;
  assign new_n2554 = \V14(0)  & new_n2553;
  assign new_n2555 = ~\V260(0)  & ~new_n2552;
  assign new_n2556 = \V14(0)  & new_n2555;
  assign \V1467(0)  = new_n2554 | new_n2556;
  assign new_n2558 = \V14(0)  & ~new_n1503;
  assign new_n2559 = new_n2254 & new_n2558;
  assign V1470 = \V67(0)  & new_n2559;
  assign new_n2561 = \V802(0)  & \V1757(0) ;
  assign new_n2562 = new_n544 & new_n2561;
  assign new_n2563 = ~new_n544 & \V1757(0) ;
  assign new_n2564 = ~new_n1584 & ~new_n2562;
  assign \V1480(0)  = new_n2563 | ~new_n2564;
  assign new_n2566 = ~\V214(0)  & \V216(0) ;
  assign new_n2567 = ~\V70(0)  & ~\V68(0) ;
  assign new_n2568 = ~\V66(0)  & new_n2567;
  assign new_n2569 = ~\V69(0)  & new_n2568;
  assign new_n2570 = \V215(0)  & \V14(0) ;
  assign new_n2571 = ~new_n2569 & new_n2570;
  assign new_n2572 = new_n2233 & new_n2571;
  assign \V1492(0)  = new_n2566 | new_n2572;
  assign new_n2574 = \V56(0)  & ~new_n545;
  assign new_n2575 = \V171(0)  & new_n2574;
  assign new_n2576 = \V278(0)  & ~new_n567;
  assign new_n2577 = ~new_n2575 & ~new_n2576;
  assign new_n2578 = \V177(0)  & new_n2577;
  assign new_n2579 = ~\V248(0)  & new_n2578;
  assign new_n2580 = ~new_n1585 & new_n2579;
  assign new_n2581 = ~\V271(0)  & ~\V274(0) ;
  assign new_n2582 = ~\V172(0)  & new_n1470;
  assign new_n2583 = ~new_n1646 & ~new_n2580;
  assign new_n2584 = ~new_n2581 & new_n2583;
  assign new_n2585 = ~new_n2582 & new_n2584;
  assign new_n2586 = new_n544 & new_n1586;
  assign new_n2587 = \V56(0)  & new_n544;
  assign new_n2588 = \V149(7)  & new_n2587;
  assign new_n2589 = ~new_n2586 & ~new_n2588;
  assign new_n2590 = new_n2251 & ~new_n2585;
  assign \V1536(0)  = ~new_n2589 | ~new_n2590;
  assign new_n2592 = new_n2251 & \V1536(0) ;
  assign new_n2593 = ~new_n1252 & ~new_n1269;
  assign new_n2594 = ~new_n1235 & new_n2593;
  assign new_n2595 = ~new_n1218 & new_n2594;
  assign new_n2596 = ~new_n1097 & new_n2595;
  assign new_n2597 = ~new_n1114 & new_n2596;
  assign new_n2598 = ~new_n1131 & new_n2597;
  assign new_n2599 = ~new_n1148 & new_n2598;
  assign new_n2600 = ~\V1536(0)  & ~new_n2599;
  assign \V1512(3)  = new_n2592 | new_n2600;
  assign new_n2602 = new_n2251 & ~new_n2261;
  assign new_n2603 = ~new_n2589 & new_n2602;
  assign new_n2604 = \V1536(0)  & ~new_n2603;
  assign new_n2605 = ~new_n1173 & ~new_n1269;
  assign new_n2606 = ~new_n1235 & new_n2605;
  assign new_n2607 = ~new_n1207 & new_n2606;
  assign new_n2608 = ~new_n1086 & new_n2607;
  assign new_n2609 = ~new_n1114 & new_n2608;
  assign new_n2610 = ~new_n916 & new_n2609;
  assign new_n2611 = ~new_n1148 & new_n2610;
  assign new_n2612 = ~\V1536(0)  & ~new_n2611;
  assign \V1512(2)  = new_n2604 | new_n2612;
  assign new_n2614 = new_n2251 & new_n2261;
  assign new_n2615 = \V1536(0)  & ~new_n2614;
  assign new_n2616 = ~new_n1252 & new_n2605;
  assign new_n2617 = ~new_n1190 & new_n2616;
  assign new_n2618 = ~new_n1001 & new_n2617;
  assign new_n2619 = ~new_n1131 & new_n2618;
  assign new_n2620 = ~new_n916 & new_n2619;
  assign new_n2621 = ~new_n1148 & new_n2620;
  assign new_n2622 = ~\V1536(0)  & ~new_n2621;
  assign \V1512(1)  = new_n2615 | new_n2622;
  assign new_n2624 = \V68(0)  & new_n2254;
  assign V1537 = \V14(0)  & new_n2624;
  assign new_n2626 = ~\V69(0)  & ~\V50(0) ;
  assign new_n2627 = new_n2254 & ~new_n2626;
  assign V1539 = \V14(0)  & new_n2627;
  assign new_n2629 = ~\V239(4)  & ~\V802(0) ;
  assign new_n2630 = new_n591 & new_n2629;
  assign new_n2631 = ~new_n2498 & new_n2630;
  assign new_n2632 = ~\V802(0)  & new_n591;
  assign new_n2633 = \V1243(9)  & ~new_n2632;
  assign new_n2634 = new_n2498 & new_n2633;
  assign \V1552(1)  = new_n2631 | new_n2634;
  assign new_n2636 = \V239(4)  & ~\V239(3) ;
  assign new_n2637 = ~\V239(4)  & \V239(3) ;
  assign new_n2638 = ~new_n2636 & ~new_n2637;
  assign new_n2639 = ~\V802(0)  & ~new_n2638;
  assign new_n2640 = new_n591 & new_n2639;
  assign new_n2641 = ~new_n2498 & new_n2640;
  assign new_n2642 = \V1243(8)  & ~new_n2632;
  assign new_n2643 = new_n2498 & new_n2642;
  assign \V1552(0)  = new_n2641 | new_n2643;
  assign new_n2645 = \V132(1)  & new_n2301;
  assign new_n2646 = ~new_n2307 & new_n2645;
  assign \V1953(1)  = ~new_n2278 & new_n2646;
  assign new_n2648 = \V132(0)  & new_n2301;
  assign new_n2649 = ~new_n2307 & new_n2648;
  assign new_n2650 = ~new_n2278 & new_n2649;
  assign new_n2651 = \V108(5)  & ~new_n2301;
  assign new_n2652 = ~new_n2307 & new_n2651;
  assign new_n2653 = new_n2278 & new_n2652;
  assign \V1953(0)  = new_n2650 | new_n2653;
  assign new_n2655 = \V1953(1)  & ~\V1953(0) ;
  assign new_n2656 = ~\V1953(1)  & \V1953(0) ;
  assign new_n2657 = ~new_n2655 & ~new_n2656;
  assign new_n2658 = \V100(5)  & new_n2306;
  assign new_n2659 = ~new_n2308 & new_n2658;
  assign new_n2660 = ~new_n2301 & new_n2659;
  assign new_n2661 = ~new_n2277 & new_n2660;
  assign new_n2662 = \V213(5)  & ~new_n2306;
  assign new_n2663 = new_n2308 & new_n2662;
  assign new_n2664 = ~new_n2301 & new_n2663;
  assign new_n2665 = ~new_n2277 & new_n2664;
  assign new_n2666 = \V124(5)  & ~new_n2306;
  assign new_n2667 = ~new_n2308 & new_n2666;
  assign new_n2668 = new_n2301 & new_n2667;
  assign new_n2669 = ~new_n2277 & new_n2668;
  assign new_n2670 = ~new_n2661 & ~new_n2665;
  assign \V1921(5)  = new_n2669 | ~new_n2670;
  assign new_n2672 = \V100(4)  & new_n2306;
  assign new_n2673 = ~new_n2308 & new_n2672;
  assign new_n2674 = ~new_n2301 & new_n2673;
  assign new_n2675 = ~new_n2277 & new_n2674;
  assign new_n2676 = \V213(4)  & ~new_n2306;
  assign new_n2677 = new_n2308 & new_n2676;
  assign new_n2678 = ~new_n2301 & new_n2677;
  assign new_n2679 = ~new_n2277 & new_n2678;
  assign new_n2680 = \V124(4)  & ~new_n2306;
  assign new_n2681 = ~new_n2308 & new_n2680;
  assign new_n2682 = new_n2301 & new_n2681;
  assign new_n2683 = ~new_n2277 & new_n2682;
  assign new_n2684 = \V108(4)  & ~new_n2306;
  assign new_n2685 = ~new_n2308 & new_n2684;
  assign new_n2686 = ~new_n2301 & new_n2685;
  assign new_n2687 = new_n2277 & new_n2686;
  assign new_n2688 = ~new_n2683 & ~new_n2687;
  assign new_n2689 = ~new_n2675 & ~new_n2679;
  assign \V1921(4)  = ~new_n2688 | ~new_n2689;
  assign new_n2691 = \V1921(5)  & ~\V1921(4) ;
  assign new_n2692 = ~\V1921(5)  & \V1921(4) ;
  assign new_n2693 = ~new_n2691 & ~new_n2692;
  assign new_n2694 = ~new_n2657 & new_n2693;
  assign new_n2695 = new_n2657 & ~new_n2693;
  assign new_n2696 = ~new_n2694 & ~new_n2695;
  assign new_n2697 = \V100(3)  & new_n2306;
  assign new_n2698 = ~new_n2308 & new_n2697;
  assign new_n2699 = ~new_n2301 & new_n2698;
  assign new_n2700 = ~new_n2277 & new_n2699;
  assign new_n2701 = \V213(3)  & ~new_n2306;
  assign new_n2702 = new_n2308 & new_n2701;
  assign new_n2703 = ~new_n2301 & new_n2702;
  assign new_n2704 = ~new_n2277 & new_n2703;
  assign new_n2705 = \V124(3)  & ~new_n2306;
  assign new_n2706 = ~new_n2308 & new_n2705;
  assign new_n2707 = new_n2301 & new_n2706;
  assign new_n2708 = ~new_n2277 & new_n2707;
  assign new_n2709 = \V108(3)  & ~new_n2306;
  assign new_n2710 = ~new_n2308 & new_n2709;
  assign new_n2711 = ~new_n2301 & new_n2710;
  assign new_n2712 = new_n2277 & new_n2711;
  assign new_n2713 = ~new_n2708 & ~new_n2712;
  assign new_n2714 = ~new_n2700 & ~new_n2704;
  assign \V1921(3)  = ~new_n2713 | ~new_n2714;
  assign new_n2716 = \V100(2)  & new_n2306;
  assign new_n2717 = ~new_n2308 & new_n2716;
  assign new_n2718 = ~new_n2301 & new_n2717;
  assign new_n2719 = ~new_n2277 & new_n2718;
  assign new_n2720 = \V213(2)  & ~new_n2306;
  assign new_n2721 = new_n2308 & new_n2720;
  assign new_n2722 = ~new_n2301 & new_n2721;
  assign new_n2723 = ~new_n2277 & new_n2722;
  assign new_n2724 = \V124(2)  & ~new_n2306;
  assign new_n2725 = ~new_n2308 & new_n2724;
  assign new_n2726 = new_n2301 & new_n2725;
  assign new_n2727 = ~new_n2277 & new_n2726;
  assign new_n2728 = \V108(2)  & ~new_n2306;
  assign new_n2729 = ~new_n2308 & new_n2728;
  assign new_n2730 = ~new_n2301 & new_n2729;
  assign new_n2731 = new_n2277 & new_n2730;
  assign new_n2732 = ~new_n2727 & ~new_n2731;
  assign new_n2733 = ~new_n2719 & ~new_n2723;
  assign \V1921(2)  = ~new_n2732 | ~new_n2733;
  assign new_n2735 = \V1921(3)  & ~\V1921(2) ;
  assign new_n2736 = ~\V1921(3)  & \V1921(2) ;
  assign new_n2737 = ~new_n2735 & ~new_n2736;
  assign new_n2738 = \V100(1)  & new_n2306;
  assign new_n2739 = ~new_n2308 & new_n2738;
  assign new_n2740 = ~new_n2301 & new_n2739;
  assign new_n2741 = ~new_n2277 & new_n2740;
  assign new_n2742 = \V213(1)  & ~new_n2306;
  assign new_n2743 = new_n2308 & new_n2742;
  assign new_n2744 = ~new_n2301 & new_n2743;
  assign new_n2745 = ~new_n2277 & new_n2744;
  assign new_n2746 = \V124(1)  & ~new_n2306;
  assign new_n2747 = ~new_n2308 & new_n2746;
  assign new_n2748 = new_n2301 & new_n2747;
  assign new_n2749 = ~new_n2277 & new_n2748;
  assign new_n2750 = \V108(1)  & ~new_n2306;
  assign new_n2751 = ~new_n2308 & new_n2750;
  assign new_n2752 = ~new_n2301 & new_n2751;
  assign new_n2753 = new_n2277 & new_n2752;
  assign new_n2754 = ~new_n2749 & ~new_n2753;
  assign new_n2755 = ~new_n2741 & ~new_n2745;
  assign \V1921(1)  = ~new_n2754 | ~new_n2755;
  assign new_n2757 = \V100(0)  & new_n2306;
  assign new_n2758 = ~new_n2308 & new_n2757;
  assign new_n2759 = ~new_n2301 & new_n2758;
  assign new_n2760 = ~new_n2277 & new_n2759;
  assign new_n2761 = \V213(0)  & ~new_n2306;
  assign new_n2762 = new_n2308 & new_n2761;
  assign new_n2763 = ~new_n2301 & new_n2762;
  assign new_n2764 = ~new_n2277 & new_n2763;
  assign new_n2765 = \V124(0)  & ~new_n2306;
  assign new_n2766 = ~new_n2308 & new_n2765;
  assign new_n2767 = new_n2301 & new_n2766;
  assign new_n2768 = ~new_n2277 & new_n2767;
  assign new_n2769 = \V108(0)  & ~new_n2306;
  assign new_n2770 = ~new_n2308 & new_n2769;
  assign new_n2771 = ~new_n2301 & new_n2770;
  assign new_n2772 = new_n2277 & new_n2771;
  assign new_n2773 = ~new_n2768 & ~new_n2772;
  assign new_n2774 = ~new_n2760 & ~new_n2764;
  assign \V1921(0)  = ~new_n2773 | ~new_n2774;
  assign new_n2776 = \V1921(1)  & ~\V1921(0) ;
  assign new_n2777 = ~\V1921(1)  & \V1921(0) ;
  assign new_n2778 = ~new_n2776 & ~new_n2777;
  assign new_n2779 = ~new_n2737 & new_n2778;
  assign new_n2780 = new_n2737 & ~new_n2778;
  assign new_n2781 = ~new_n2779 & ~new_n2780;
  assign new_n2782 = ~new_n2696 & new_n2781;
  assign new_n2783 = new_n2696 & ~new_n2781;
  assign \V1613(0)  = ~new_n2782 & ~new_n2783;
  assign new_n2785 = \V118(7)  & new_n2307;
  assign new_n2786 = new_n1628 & new_n2785;
  assign new_n2787 = \V46(0)  & ~new_n2307;
  assign new_n2788 = ~new_n1628 & new_n2787;
  assign \V1960(1)  = new_n2786 | new_n2788;
  assign new_n2790 = \V118(6)  & new_n2307;
  assign new_n2791 = new_n1628 & new_n2790;
  assign new_n2792 = \V48(0)  & ~new_n2307;
  assign new_n2793 = ~new_n1628 & new_n2792;
  assign \V1960(0)  = new_n2791 | new_n2793;
  assign new_n2795 = \V1960(1)  & ~\V1960(0) ;
  assign new_n2796 = ~\V1960(1)  & \V1960(0) ;
  assign new_n2797 = ~new_n2795 & ~new_n2796;
  assign new_n2798 = \V132(7)  & new_n2301;
  assign new_n2799 = ~new_n2307 & new_n2798;
  assign new_n2800 = ~new_n2278 & new_n2799;
  assign new_n2801 = \V118(5)  & ~new_n2301;
  assign new_n2802 = new_n2307 & new_n2801;
  assign new_n2803 = ~new_n2278 & new_n2802;
  assign \V1953(7)  = new_n2800 | new_n2803;
  assign new_n2805 = \V132(6)  & new_n2301;
  assign new_n2806 = ~new_n2307 & new_n2805;
  assign new_n2807 = ~new_n2278 & new_n2806;
  assign new_n2808 = \V118(4)  & ~new_n2301;
  assign new_n2809 = new_n2307 & new_n2808;
  assign new_n2810 = ~new_n2278 & new_n2809;
  assign \V1953(6)  = new_n2807 | new_n2810;
  assign new_n2812 = \V1953(7)  & ~\V1953(6) ;
  assign new_n2813 = ~\V1953(7)  & \V1953(6) ;
  assign new_n2814 = ~new_n2812 & ~new_n2813;
  assign new_n2815 = ~new_n2797 & new_n2814;
  assign new_n2816 = new_n2797 & ~new_n2814;
  assign new_n2817 = ~new_n2815 & ~new_n2816;
  assign new_n2818 = \V132(5)  & new_n2301;
  assign new_n2819 = ~new_n2307 & new_n2818;
  assign new_n2820 = ~new_n2278 & new_n2819;
  assign new_n2821 = \V118(3)  & ~new_n2301;
  assign new_n2822 = new_n2307 & new_n2821;
  assign new_n2823 = ~new_n2278 & new_n2822;
  assign \V1953(5)  = new_n2820 | new_n2823;
  assign new_n2825 = \V132(4)  & new_n2301;
  assign new_n2826 = ~new_n2307 & new_n2825;
  assign new_n2827 = ~new_n2278 & new_n2826;
  assign new_n2828 = \V118(2)  & ~new_n2301;
  assign new_n2829 = new_n2307 & new_n2828;
  assign new_n2830 = ~new_n2278 & new_n2829;
  assign \V1953(4)  = new_n2827 | new_n2830;
  assign new_n2832 = \V1953(5)  & ~\V1953(4) ;
  assign new_n2833 = ~\V1953(5)  & \V1953(4) ;
  assign new_n2834 = ~new_n2832 & ~new_n2833;
  assign new_n2835 = \V132(3)  & new_n2301;
  assign new_n2836 = ~new_n2307 & new_n2835;
  assign new_n2837 = ~new_n2278 & new_n2836;
  assign new_n2838 = \V118(1)  & ~new_n2301;
  assign new_n2839 = new_n2307 & new_n2838;
  assign new_n2840 = ~new_n2278 & new_n2839;
  assign \V1953(3)  = new_n2837 | new_n2840;
  assign new_n2842 = \V132(2)  & new_n2301;
  assign new_n2843 = ~new_n2307 & new_n2842;
  assign new_n2844 = ~new_n2278 & new_n2843;
  assign new_n2845 = \V118(0)  & ~new_n2301;
  assign new_n2846 = new_n2307 & new_n2845;
  assign new_n2847 = ~new_n2278 & new_n2846;
  assign \V1953(2)  = new_n2844 | new_n2847;
  assign new_n2849 = \V1953(3)  & ~\V1953(2) ;
  assign new_n2850 = ~\V1953(3)  & \V1953(2) ;
  assign new_n2851 = ~new_n2849 & ~new_n2850;
  assign new_n2852 = ~new_n2834 & new_n2851;
  assign new_n2853 = new_n2834 & ~new_n2851;
  assign new_n2854 = ~new_n2852 & ~new_n2853;
  assign new_n2855 = ~new_n2817 & new_n2854;
  assign new_n2856 = new_n2817 & ~new_n2854;
  assign \V1613(1)  = ~new_n2855 & ~new_n2856;
  assign new_n2858 = \V174(0)  & new_n1311;
  assign new_n2859 = ~\V302(0)  & \V292(0) ;
  assign new_n2860 = \V174(0)  & ~new_n2251;
  assign new_n2861 = ~new_n2859 & ~new_n2860;
  assign new_n2862 = ~new_n509 & ~new_n2858;
  assign \V1620(0)  = ~new_n2861 | ~new_n2862;
  assign new_n2864 = \V62(0)  & \V91(1) ;
  assign new_n2865 = \V59(0)  & \V91(0) ;
  assign new_n2866 = ~new_n2864 & ~new_n2865;
  assign new_n2867 = new_n1514 & ~new_n2866;
  assign new_n2868 = ~\V294(0)  & ~new_n1513;
  assign new_n2869 = ~new_n1620 & new_n2868;
  assign new_n2870 = new_n2197 & ~new_n2867;
  assign \V1629(0)  = new_n2869 | ~new_n2870;
  assign new_n2872 = \V149(7)  & new_n1508;
  assign new_n2873 = ~new_n2424 & ~new_n2872;
  assign \V1645(0)  = new_n1523 | ~new_n2873;
  assign new_n2875 = ~\V289(0)  & new_n534;
  assign new_n2876 = ~\V249(0)  & new_n2875;
  assign new_n2877 = ~new_n1609 & new_n2876;
  assign new_n2878 = \V295(0)  & new_n2877;
  assign \V1652(0)  = \V290(0)  | ~new_n2878;
  assign new_n2880 = ~\V59(0)  & ~\V259(0) ;
  assign new_n2881 = ~\V260(0)  & new_n2880;
  assign new_n2882 = \V258(0)  & new_n2881;
  assign new_n2883 = \V14(0)  & \V262(0) ;
  assign new_n2884 = ~new_n2882 & new_n2883;
  assign new_n2885 = \V262(0)  & new_n2884;
  assign new_n2886 = new_n533 & ~new_n2885;
  assign new_n2887 = ~new_n2301 & ~new_n2308;
  assign new_n2888 = ~new_n1576 & new_n2886;
  assign new_n2889 = new_n2887 & new_n2888;
  assign new_n2890 = ~new_n2306 & ~new_n2307;
  assign new_n2891 = ~new_n2300 & new_n2890;
  assign new_n2892 = new_n2889 & new_n2891;
  assign new_n2893 = ~\V289(0)  & new_n2892;
  assign new_n2894 = \V1741(0)  & new_n2893;
  assign new_n2895 = new_n2317 & new_n2892;
  assign new_n2896 = new_n2886 & new_n2895;
  assign new_n2897 = ~new_n1513 & new_n2896;
  assign new_n2898 = ~\V289(0)  & new_n2320;
  assign new_n2899 = new_n2251 & new_n2898;
  assign new_n2900 = ~new_n2897 & new_n2899;
  assign new_n2901 = ~new_n2207 & new_n2900;
  assign new_n2902 = ~\V289(0)  & new_n1457;
  assign new_n2903 = ~\V802(0)  & new_n2902;
  assign new_n2904 = ~new_n1504 & ~new_n2894;
  assign new_n2905 = ~new_n2901 & new_n2904;
  assign V1669 = ~new_n2903 & new_n2905;
  assign \V1679(0)  = ~new_n533 | new_n2884;
  assign new_n2908 = \V56(0)  & new_n2306;
  assign new_n2909 = ~new_n487 & ~new_n489;
  assign new_n2910 = new_n1311 & ~new_n2909;
  assign new_n2911 = \V290(0)  & new_n2910;
  assign new_n2912 = ~new_n1311 & ~new_n2909;
  assign new_n2913 = new_n1586 & new_n2912;
  assign new_n2914 = ~new_n2424 & new_n2913;
  assign new_n2915 = ~new_n499 & new_n2914;
  assign new_n2916 = ~new_n2911 & ~new_n2915;
  assign new_n2917 = \V14(0)  & ~new_n2908;
  assign new_n2918 = \V100(0)  & new_n2917;
  assign new_n2919 = new_n2916 & new_n2918;
  assign new_n2920 = new_n2916 & new_n2919;
  assign new_n2921 = ~new_n2439 & ~new_n2916;
  assign new_n2922 = ~new_n2916 & new_n2921;
  assign \V1693(0)  = new_n2920 | new_n2922;
  assign new_n2924 = \V100(5)  & new_n2917;
  assign new_n2925 = ~new_n2911 & new_n2924;
  assign new_n2926 = ~new_n2911 & new_n2925;
  assign new_n2927 = \V165(7)  & new_n2911;
  assign new_n2928 = new_n2911 & new_n2927;
  assign \V1709(4)  = new_n2926 | new_n2928;
  assign new_n2930 = \V100(4)  & new_n2917;
  assign new_n2931 = ~new_n2911 & new_n2930;
  assign new_n2932 = ~new_n2911 & new_n2931;
  assign new_n2933 = \V165(6)  & new_n2911;
  assign new_n2934 = new_n2911 & new_n2933;
  assign \V1709(3)  = new_n2932 | new_n2934;
  assign new_n2936 = \V100(3)  & new_n2917;
  assign new_n2937 = ~new_n2911 & new_n2936;
  assign new_n2938 = ~new_n2911 & new_n2937;
  assign new_n2939 = \V165(5)  & new_n2911;
  assign new_n2940 = new_n2911 & new_n2939;
  assign \V1709(2)  = new_n2938 | new_n2940;
  assign new_n2942 = \V100(2)  & new_n2917;
  assign new_n2943 = ~new_n2911 & new_n2942;
  assign new_n2944 = ~new_n2911 & new_n2943;
  assign new_n2945 = \V165(4)  & new_n2911;
  assign new_n2946 = new_n2911 & new_n2945;
  assign \V1709(1)  = new_n2944 | new_n2946;
  assign new_n2948 = \V100(1)  & new_n2917;
  assign new_n2949 = ~new_n2911 & new_n2948;
  assign new_n2950 = ~new_n2911 & new_n2949;
  assign new_n2951 = \V165(3)  & new_n2911;
  assign new_n2952 = new_n2911 & new_n2951;
  assign \V1709(0)  = new_n2950 | new_n2952;
  assign new_n2954 = ~\V280(0)  & new_n591;
  assign new_n2955 = ~new_n1304 & ~new_n1311;
  assign new_n2956 = new_n2254 & new_n2955;
  assign new_n2957 = ~new_n2954 & new_n2956;
  assign new_n2958 = \V240(0)  & new_n2957;
  assign new_n2959 = ~\V172(0)  & new_n2958;
  assign new_n2960 = ~new_n591 & ~new_n1421;
  assign new_n2961 = \V802(0)  & ~new_n2960;
  assign \V1717(0)  = new_n2959 | new_n2961;
  assign new_n2963 = \V14(0)  & \V242(0) ;
  assign new_n2964 = new_n566 & new_n2963;
  assign new_n2965 = ~new_n567 & new_n1858;
  assign new_n2966 = ~\V1536(0)  & new_n2965;
  assign \V1726(0)  = new_n2964 | new_n2966;
  assign new_n2968 = new_n1604 & new_n2902;
  assign new_n2969 = ~\V802(0)  & new_n2968;
  assign V1736 = ~\V290(0)  & new_n2969;
  assign new_n2971 = \V33(0)  & ~new_n499;
  assign new_n2972 = \V289(0)  & new_n2971;
  assign \V1745(0)  = new_n485 | ~new_n2972;
  assign new_n2974 = \V16(0)  & ~\V15(0) ;
  assign \V1758(0)  = new_n1474 | new_n2974;
  assign new_n2976 = new_n485 & new_n2974;
  assign new_n2977 = new_n487 & new_n2974;
  assign new_n2978 = \V56(0)  & new_n2278;
  assign new_n2979 = \V101(0)  & ~new_n2978;
  assign new_n2980 = \V14(0)  & new_n2979;
  assign new_n2981 = ~new_n2976 & ~new_n2977;
  assign \V1759(0)  = new_n2980 | ~new_n2981;
  assign new_n2983 = ~\V88(3)  & new_n598;
  assign new_n2984 = new_n598 & new_n2983;
  assign new_n2985 = ~\V134(1)  & ~new_n598;
  assign new_n2986 = ~new_n598 & new_n2985;
  assign \V1771(1)  = new_n2984 | new_n2986;
  assign new_n2988 = ~\V88(2)  & new_n598;
  assign new_n2989 = new_n598 & new_n2988;
  assign new_n2990 = ~\V134(0)  & ~new_n598;
  assign new_n2991 = ~new_n598 & new_n2990;
  assign \V1771(0)  = new_n2989 | new_n2991;
  assign new_n2993 = ~new_n598 & ~\V1213(11) ;
  assign new_n2994 = ~new_n598 & new_n2993;
  assign new_n2995 = ~\V78(3)  & new_n598;
  assign new_n2996 = new_n598 & new_n2995;
  assign \V1781(1)  = new_n2994 | new_n2996;
  assign new_n2998 = ~new_n598 & ~\V1213(10) ;
  assign new_n2999 = ~new_n598 & new_n2998;
  assign new_n3000 = ~\V78(2)  & new_n598;
  assign new_n3001 = new_n598 & new_n3000;
  assign \V1781(0)  = new_n2999 | new_n3001;
  assign new_n3003 = \V37(0)  & ~\V1243(9) ;
  assign new_n3004 = \V37(0)  & new_n3003;
  assign new_n3005 = ~\V37(0)  & \V321(2) ;
  assign new_n3006 = ~\V37(0)  & new_n3005;
  assign \V1829(9)  = new_n3004 | new_n3006;
  assign new_n3008 = \V37(0)  & ~\V1243(8) ;
  assign new_n3009 = \V37(0)  & new_n3008;
  assign new_n3010 = ~\V37(0)  & ~\V1213(11) ;
  assign new_n3011 = ~\V37(0)  & new_n3010;
  assign \V1829(8)  = new_n3009 | new_n3011;
  assign new_n3013 = \V37(0)  & ~\V1243(7) ;
  assign new_n3014 = \V37(0)  & new_n3013;
  assign new_n3015 = ~\V37(0)  & ~\V1213(10) ;
  assign new_n3016 = ~\V37(0)  & new_n3015;
  assign \V1829(7)  = new_n3014 | new_n3016;
  assign new_n3018 = \V37(0)  & ~\V1243(6) ;
  assign new_n3019 = \V37(0)  & new_n3018;
  assign new_n3020 = ~\V37(0)  & ~\V1213(9) ;
  assign new_n3021 = ~\V37(0)  & new_n3020;
  assign \V1829(6)  = new_n3019 | new_n3021;
  assign new_n3023 = \V37(0)  & ~\V1243(5) ;
  assign new_n3024 = \V37(0)  & new_n3023;
  assign new_n3025 = ~\V37(0)  & ~\V1213(8) ;
  assign new_n3026 = ~\V37(0)  & new_n3025;
  assign \V1829(5)  = new_n3024 | new_n3026;
  assign new_n3028 = \V37(0)  & ~\V1243(4) ;
  assign new_n3029 = \V37(0)  & new_n3028;
  assign new_n3030 = ~\V37(0)  & ~\V1213(7) ;
  assign new_n3031 = ~\V37(0)  & new_n3030;
  assign \V1829(4)  = new_n3029 | new_n3031;
  assign new_n3033 = \V37(0)  & ~\V1243(3) ;
  assign new_n3034 = \V37(0)  & new_n3033;
  assign new_n3035 = ~\V37(0)  & ~\V1213(6) ;
  assign new_n3036 = ~\V37(0)  & new_n3035;
  assign \V1829(3)  = new_n3034 | new_n3036;
  assign new_n3038 = \V37(0)  & ~\V1243(2) ;
  assign new_n3039 = \V37(0)  & new_n3038;
  assign new_n3040 = ~\V37(0)  & ~\V1213(5) ;
  assign new_n3041 = ~\V37(0)  & new_n3040;
  assign \V1829(2)  = new_n3039 | new_n3041;
  assign new_n3043 = \V37(0)  & ~\V1243(1) ;
  assign new_n3044 = \V37(0)  & new_n3043;
  assign new_n3045 = ~\V37(0)  & ~\V1213(4) ;
  assign new_n3046 = ~\V37(0)  & new_n3045;
  assign \V1829(1)  = new_n3044 | new_n3046;
  assign new_n3048 = \V37(0)  & ~\V1213(2) ;
  assign new_n3049 = \V37(0)  & new_n3048;
  assign \V1829(0)  = new_n3006 | new_n3049;
  assign new_n3051 = \V262(0)  & ~new_n2884;
  assign new_n3052 = ~new_n2508 & new_n3051;
  assign new_n3053 = \V261(0)  & ~new_n3052;
  assign new_n3054 = ~new_n2535 & ~new_n3053;
  assign V1832 = \V14(0)  & ~new_n3054;
  assign new_n3056 = \V56(0)  & new_n2277;
  assign new_n3057 = \V108(0)  & ~new_n3056;
  assign new_n3058 = ~new_n1584 & ~new_n3057;
  assign \V1896(0)  = new_n1475 | ~new_n3058;
  assign new_n3060 = new_n538 & new_n1584;
  assign new_n3061 = \V108(1)  & ~new_n3056;
  assign \V1897(0)  = new_n3060 | new_n3061;
  assign new_n3063 = new_n485 & new_n2221;
  assign new_n3064 = \V108(2)  & ~new_n3056;
  assign \V1898(0)  = new_n3063 | new_n3064;
  assign new_n3066 = new_n487 & new_n2221;
  assign new_n3067 = \V108(3)  & ~new_n3056;
  assign \V1899(0)  = new_n3066 | new_n3067;
  assign new_n3069 = \V108(4)  & ~new_n3056;
  assign \V1900(0)  = new_n1474 | new_n3069;
  assign new_n3071 = \V108(5)  & ~new_n2978;
  assign \V1901(0)  = new_n2974 | new_n3071;
  assign new_n3073 = ~\V108(4)  & new_n1474;
  assign new_n3074 = \V101(0)  & new_n3073;
  assign new_n3075 = \V56(0)  & new_n2307;
  assign new_n3076 = \V110(0)  & ~new_n3074;
  assign new_n3077 = ~new_n3075 & new_n3076;
  assign new_n3078 = \V14(0)  & new_n3077;
  assign new_n3079 = ~\V102(0)  & ~\V1758(0) ;
  assign new_n3080 = ~\V110(0)  & ~new_n3079;
  assign new_n3081 = new_n487 & new_n3080;
  assign \V1968(0)  = new_n3078 | new_n3081;
  assign new_n3083 = ~new_n1860 & ~new_n2481;
  assign new_n3084 = ~\V134(1)  & ~new_n2481;
  assign new_n3085 = new_n1860 & new_n3084;
  assign new_n3086 = ~new_n3083 & new_n3085;
  assign new_n3087 = new_n1860 & ~new_n2481;
  assign new_n3088 = \V134(1)  & ~new_n1860;
  assign new_n3089 = ~new_n2481 & new_n3088;
  assign new_n3090 = ~new_n3087 & new_n3089;
  assign \V1992(1)  = new_n3086 | new_n3090;
  assign new_n3092 = \V134(1)  & ~\V134(0) ;
  assign new_n3093 = ~\V134(1)  & \V134(0) ;
  assign new_n3094 = ~new_n3092 & ~new_n3093;
  assign new_n3095 = ~new_n2481 & ~new_n3094;
  assign new_n3096 = new_n1860 & new_n3095;
  assign new_n3097 = ~new_n3083 & new_n3096;
  assign new_n3098 = \V134(0)  & ~new_n1860;
  assign new_n3099 = ~new_n2481 & new_n3098;
  assign new_n3100 = ~new_n3087 & new_n3099;
  assign \V1992(0)  = new_n3097 | new_n3100;
  assign new_n3102 = \V257(7)  & \V257(5) ;
  assign new_n3103 = \V257(3)  & new_n3102;
  assign new_n3104 = \V257(1)  & new_n3103;
  assign new_n3105 = \V257(2)  & new_n3104;
  assign new_n3106 = \V257(4)  & new_n3105;
  assign new_n3107 = \V257(6)  & new_n3106;
  assign new_n3108 = \V257(0)  & ~new_n3107;
  assign new_n3109 = ~\V257(0)  & new_n3107;
  assign V650 = new_n3108 | new_n3109;
  assign new_n3111 = \V257(2)  & new_n3103;
  assign new_n3112 = \V257(4)  & new_n3111;
  assign new_n3113 = \V257(6)  & new_n3112;
  assign new_n3114 = \V257(1)  & ~new_n3113;
  assign new_n3115 = ~\V257(1)  & new_n3113;
  assign V651 = new_n3114 | new_n3115;
  assign new_n3117 = \V257(4)  & new_n3103;
  assign new_n3118 = \V257(6)  & new_n3117;
  assign new_n3119 = \V257(2)  & ~new_n3118;
  assign new_n3120 = ~\V257(2)  & new_n3118;
  assign V652 = new_n3119 | new_n3120;
  assign new_n3122 = \V257(4)  & new_n3102;
  assign new_n3123 = \V257(6)  & new_n3122;
  assign new_n3124 = \V257(3)  & ~new_n3123;
  assign new_n3125 = ~\V257(3)  & new_n3123;
  assign V653 = new_n3124 | new_n3125;
  assign new_n3127 = \V257(6)  & new_n3102;
  assign new_n3128 = \V257(4)  & ~new_n3127;
  assign new_n3129 = ~\V257(4)  & new_n3127;
  assign V654 = new_n3128 | new_n3129;
  assign new_n3131 = \V257(7)  & \V257(6) ;
  assign new_n3132 = \V257(5)  & ~new_n3131;
  assign new_n3133 = ~\V257(5)  & new_n3131;
  assign V655 = new_n3132 | new_n3133;
  assign new_n3135 = ~\V257(7)  & \V257(6) ;
  assign new_n3136 = \V257(7)  & ~\V257(6) ;
  assign V656 = new_n3135 | new_n3136;
  assign new_n3138 = \V268(0)  & ~new_n2534;
  assign new_n3139 = ~\V268(0)  & new_n2534;
  assign V1370 = new_n3138 | new_n3139;
  assign new_n3141 = \V268(2)  & new_n2531;
  assign new_n3142 = \V268(4)  & new_n3141;
  assign new_n3143 = \V268(1)  & ~new_n3142;
  assign new_n3144 = ~\V268(1)  & new_n3142;
  assign V1371 = new_n3143 | new_n3144;
  assign new_n3146 = \V268(4)  & new_n2531;
  assign new_n3147 = \V268(2)  & ~new_n3146;
  assign new_n3148 = ~\V268(2)  & new_n3146;
  assign V1372 = new_n3147 | new_n3148;
  assign new_n3150 = \V268(5)  & \V268(4) ;
  assign new_n3151 = \V268(3)  & ~new_n3150;
  assign new_n3152 = ~\V268(3)  & new_n3150;
  assign V1373 = new_n3151 | new_n3152;
  assign new_n3154 = ~\V268(5)  & \V268(4) ;
  assign new_n3155 = \V268(5)  & ~\V268(4) ;
  assign V1374 = new_n3154 | new_n3155;
  assign \V585(0)  = ~\V34(0) ;
  assign V657 = ~\V257(7) ;
  assign \V1243(0)  = ~\V321(2) ;
  assign V1375 = ~\V268(5) ;
  assign \V1481(0)  = ~\V214(0) ;
  assign \V1495(0)  = ~\V175(0) ;
  assign \V1671(0)  = ~\V205(0) ;
  assign \V1760(0)  = ~\V101(0) ;
  assign \V1833(0)  = ~\V261(0) ;
  assign \V1863(0)  = ~\V301(0) ;
  assign \V1864(0)  = ~\V302(0) ;
endmodule


