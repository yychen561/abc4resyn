// Benchmark "test" written by ABC on Tue Jan 21 21:17:19 2025

module test ( 
    i1, i2, i3, i4,
    o1  );
  input  i1, i2, i3, i4;
  output o1;
  assign o1 = i4;
endmodule


